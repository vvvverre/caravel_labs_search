magic
tech sky130B
magscale 1 2
timestamp 1660399113
<< nwell >>
rect 1066 447429 448906 447750
rect 1066 446341 448906 446907
rect 1066 445253 448906 445819
rect 1066 444165 448906 444731
rect 1066 443077 448906 443643
rect 1066 441989 448906 442555
rect 1066 440901 448906 441467
rect 1066 439813 448906 440379
rect 1066 438725 448906 439291
rect 1066 437637 448906 438203
rect 1066 436549 448906 437115
rect 1066 435461 448906 436027
rect 1066 434373 448906 434939
rect 1066 433285 448906 433851
rect 1066 432197 448906 432763
rect 1066 431109 448906 431675
rect 1066 430021 448906 430587
rect 1066 428933 448906 429499
rect 1066 427845 448906 428411
rect 1066 426757 448906 427323
rect 1066 425669 448906 426235
rect 1066 424581 448906 425147
rect 1066 423493 448906 424059
rect 1066 422405 448906 422971
rect 1066 421317 448906 421883
rect 1066 420229 448906 420795
rect 1066 419141 448906 419707
rect 1066 418053 448906 418619
rect 1066 416965 448906 417531
rect 1066 415877 448906 416443
rect 1066 414789 448906 415355
rect 1066 413701 448906 414267
rect 1066 412613 448906 413179
rect 1066 411525 448906 412091
rect 1066 410437 448906 411003
rect 1066 409349 448906 409915
rect 1066 408261 448906 408827
rect 1066 407173 448906 407739
rect 1066 406085 448906 406651
rect 1066 404997 448906 405563
rect 1066 403909 448906 404475
rect 1066 402821 448906 403387
rect 1066 401733 448906 402299
rect 1066 400645 448906 401211
rect 1066 399557 448906 400123
rect 1066 398469 448906 399035
rect 1066 397381 448906 397947
rect 1066 396293 448906 396859
rect 1066 395205 448906 395771
rect 1066 394117 448906 394683
rect 1066 393029 448906 393595
rect 1066 391941 448906 392507
rect 1066 390853 448906 391419
rect 1066 389765 448906 390331
rect 1066 388677 448906 389243
rect 1066 387589 448906 388155
rect 1066 386501 448906 387067
rect 1066 385413 448906 385979
rect 1066 384325 448906 384891
rect 1066 383237 448906 383803
rect 1066 382149 448906 382715
rect 1066 381061 448906 381627
rect 1066 379973 448906 380539
rect 1066 378885 448906 379451
rect 1066 377797 448906 378363
rect 1066 376709 448906 377275
rect 1066 375621 448906 376187
rect 1066 374533 448906 375099
rect 1066 373445 448906 374011
rect 1066 372357 448906 372923
rect 1066 371269 448906 371835
rect 1066 370181 448906 370747
rect 1066 369093 448906 369659
rect 1066 368005 448906 368571
rect 1066 366917 448906 367483
rect 1066 365829 448906 366395
rect 1066 364741 448906 365307
rect 1066 363653 448906 364219
rect 1066 362565 448906 363131
rect 1066 361477 448906 362043
rect 1066 360389 448906 360955
rect 1066 359301 448906 359867
rect 1066 358213 448906 358779
rect 1066 357125 448906 357691
rect 1066 356037 448906 356603
rect 1066 354949 448906 355515
rect 1066 353861 448906 354427
rect 1066 352773 448906 353339
rect 1066 351685 448906 352251
rect 1066 350597 448906 351163
rect 1066 349509 448906 350075
rect 1066 348421 448906 348987
rect 1066 347333 448906 347899
rect 1066 346245 448906 346811
rect 1066 345157 448906 345723
rect 1066 344069 448906 344635
rect 1066 342981 448906 343547
rect 1066 341893 448906 342459
rect 1066 340805 448906 341371
rect 1066 339717 448906 340283
rect 1066 338629 448906 339195
rect 1066 337541 448906 338107
rect 1066 336453 448906 337019
rect 1066 335365 448906 335931
rect 1066 334277 448906 334843
rect 1066 333189 448906 333755
rect 1066 332101 448906 332667
rect 1066 331013 448906 331579
rect 1066 329925 448906 330491
rect 1066 328837 448906 329403
rect 1066 327749 448906 328315
rect 1066 326661 448906 327227
rect 1066 325573 448906 326139
rect 1066 324485 448906 325051
rect 1066 323397 448906 323963
rect 1066 322309 448906 322875
rect 1066 321221 448906 321787
rect 1066 320133 448906 320699
rect 1066 319045 448906 319611
rect 1066 317957 448906 318523
rect 1066 316869 448906 317435
rect 1066 315781 448906 316347
rect 1066 314693 448906 315259
rect 1066 313605 448906 314171
rect 1066 312517 448906 313083
rect 1066 311429 448906 311995
rect 1066 310341 448906 310907
rect 1066 309253 448906 309819
rect 1066 308165 448906 308731
rect 1066 307077 448906 307643
rect 1066 305989 448906 306555
rect 1066 304901 448906 305467
rect 1066 303813 448906 304379
rect 1066 302725 448906 303291
rect 1066 301637 448906 302203
rect 1066 300549 448906 301115
rect 1066 299461 448906 300027
rect 1066 298373 448906 298939
rect 1066 297285 448906 297851
rect 1066 296197 448906 296763
rect 1066 295109 448906 295675
rect 1066 294021 448906 294587
rect 1066 292933 448906 293499
rect 1066 291845 448906 292411
rect 1066 290757 448906 291323
rect 1066 289669 448906 290235
rect 1066 288581 448906 289147
rect 1066 287493 448906 288059
rect 1066 286405 448906 286971
rect 1066 285317 448906 285883
rect 1066 284229 448906 284795
rect 1066 283141 448906 283707
rect 1066 282053 448906 282619
rect 1066 280965 448906 281531
rect 1066 279877 448906 280443
rect 1066 278789 448906 279355
rect 1066 277701 448906 278267
rect 1066 276613 448906 277179
rect 1066 275525 448906 276091
rect 1066 274437 448906 275003
rect 1066 273349 448906 273915
rect 1066 272261 448906 272827
rect 1066 271173 448906 271739
rect 1066 270085 448906 270651
rect 1066 268997 448906 269563
rect 1066 267909 448906 268475
rect 1066 266821 448906 267387
rect 1066 265733 448906 266299
rect 1066 264645 448906 265211
rect 1066 263557 448906 264123
rect 1066 262469 448906 263035
rect 1066 261381 448906 261947
rect 1066 260293 448906 260859
rect 1066 259205 448906 259771
rect 1066 258117 448906 258683
rect 1066 257029 448906 257595
rect 1066 255941 448906 256507
rect 1066 254853 448906 255419
rect 1066 253765 448906 254331
rect 1066 252677 448906 253243
rect 1066 251589 448906 252155
rect 1066 250501 448906 251067
rect 1066 249413 448906 249979
rect 1066 248325 448906 248891
rect 1066 247237 448906 247803
rect 1066 246149 448906 246715
rect 1066 245061 448906 245627
rect 1066 243973 448906 244539
rect 1066 242885 448906 243451
rect 1066 241797 448906 242363
rect 1066 240709 448906 241275
rect 1066 239621 448906 240187
rect 1066 238533 448906 239099
rect 1066 237445 448906 238011
rect 1066 236357 448906 236923
rect 1066 235269 448906 235835
rect 1066 234181 448906 234747
rect 1066 233093 448906 233659
rect 1066 232005 448906 232571
rect 1066 230917 448906 231483
rect 1066 229829 448906 230395
rect 1066 228741 448906 229307
rect 1066 227653 448906 228219
rect 1066 226565 448906 227131
rect 1066 225477 448906 226043
rect 1066 224389 448906 224955
rect 1066 223301 448906 223867
rect 1066 222213 448906 222779
rect 1066 221125 448906 221691
rect 1066 220037 448906 220603
rect 1066 218949 448906 219515
rect 1066 217861 448906 218427
rect 1066 216773 448906 217339
rect 1066 215685 448906 216251
rect 1066 214597 448906 215163
rect 1066 213509 448906 214075
rect 1066 212421 448906 212987
rect 1066 211333 448906 211899
rect 1066 210245 448906 210811
rect 1066 209157 448906 209723
rect 1066 208069 448906 208635
rect 1066 206981 448906 207547
rect 1066 205893 448906 206459
rect 1066 204805 448906 205371
rect 1066 203717 448906 204283
rect 1066 202629 448906 203195
rect 1066 201541 448906 202107
rect 1066 200453 448906 201019
rect 1066 199365 448906 199931
rect 1066 198277 448906 198843
rect 1066 197189 448906 197755
rect 1066 196101 448906 196667
rect 1066 195013 448906 195579
rect 1066 193925 448906 194491
rect 1066 192837 448906 193403
rect 1066 191749 448906 192315
rect 1066 190661 448906 191227
rect 1066 189573 448906 190139
rect 1066 188485 448906 189051
rect 1066 187397 448906 187963
rect 1066 186309 448906 186875
rect 1066 185221 448906 185787
rect 1066 184133 448906 184699
rect 1066 183045 448906 183611
rect 1066 181957 448906 182523
rect 1066 180869 448906 181435
rect 1066 179781 448906 180347
rect 1066 178693 448906 179259
rect 1066 177605 448906 178171
rect 1066 176517 448906 177083
rect 1066 175429 448906 175995
rect 1066 174341 448906 174907
rect 1066 173253 448906 173819
rect 1066 172165 448906 172731
rect 1066 171077 448906 171643
rect 1066 169989 448906 170555
rect 1066 168901 448906 169467
rect 1066 167813 448906 168379
rect 1066 166725 448906 167291
rect 1066 165637 448906 166203
rect 1066 164549 448906 165115
rect 1066 163461 448906 164027
rect 1066 162373 448906 162939
rect 1066 161285 448906 161851
rect 1066 160197 448906 160763
rect 1066 159109 448906 159675
rect 1066 158021 448906 158587
rect 1066 156933 448906 157499
rect 1066 155845 448906 156411
rect 1066 154757 448906 155323
rect 1066 153669 448906 154235
rect 1066 152581 448906 153147
rect 1066 151493 448906 152059
rect 1066 150405 448906 150971
rect 1066 149317 448906 149883
rect 1066 148229 448906 148795
rect 1066 147141 448906 147707
rect 1066 146053 448906 146619
rect 1066 144965 448906 145531
rect 1066 143877 448906 144443
rect 1066 142789 448906 143355
rect 1066 141701 448906 142267
rect 1066 140613 448906 141179
rect 1066 139525 448906 140091
rect 1066 138437 448906 139003
rect 1066 137349 448906 137915
rect 1066 136261 448906 136827
rect 1066 135173 448906 135739
rect 1066 134085 448906 134651
rect 1066 132997 448906 133563
rect 1066 131909 448906 132475
rect 1066 130821 448906 131387
rect 1066 129733 448906 130299
rect 1066 128645 448906 129211
rect 1066 127557 448906 128123
rect 1066 126469 448906 127035
rect 1066 125381 448906 125947
rect 1066 124293 448906 124859
rect 1066 123205 448906 123771
rect 1066 122117 448906 122683
rect 1066 121029 448906 121595
rect 1066 119941 448906 120507
rect 1066 118853 448906 119419
rect 1066 117765 448906 118331
rect 1066 116677 448906 117243
rect 1066 115589 448906 116155
rect 1066 114501 448906 115067
rect 1066 113413 448906 113979
rect 1066 112325 448906 112891
rect 1066 111237 448906 111803
rect 1066 110149 448906 110715
rect 1066 109061 448906 109627
rect 1066 107973 448906 108539
rect 1066 106885 448906 107451
rect 1066 105797 448906 106363
rect 1066 104709 448906 105275
rect 1066 103621 448906 104187
rect 1066 102533 448906 103099
rect 1066 101445 448906 102011
rect 1066 100357 448906 100923
rect 1066 99269 448906 99835
rect 1066 98181 448906 98747
rect 1066 97093 448906 97659
rect 1066 96005 448906 96571
rect 1066 94917 448906 95483
rect 1066 93829 448906 94395
rect 1066 92741 448906 93307
rect 1066 91653 448906 92219
rect 1066 90565 448906 91131
rect 1066 89477 448906 90043
rect 1066 88389 448906 88955
rect 1066 87301 448906 87867
rect 1066 86213 448906 86779
rect 1066 85125 448906 85691
rect 1066 84037 448906 84603
rect 1066 82949 448906 83515
rect 1066 81861 448906 82427
rect 1066 80773 448906 81339
rect 1066 79685 448906 80251
rect 1066 78597 448906 79163
rect 1066 77509 448906 78075
rect 1066 76421 448906 76987
rect 1066 75333 448906 75899
rect 1066 74245 448906 74811
rect 1066 73157 448906 73723
rect 1066 72069 448906 72635
rect 1066 70981 448906 71547
rect 1066 69893 448906 70459
rect 1066 68805 448906 69371
rect 1066 67717 448906 68283
rect 1066 66629 448906 67195
rect 1066 65541 448906 66107
rect 1066 64453 448906 65019
rect 1066 63365 448906 63931
rect 1066 62277 448906 62843
rect 1066 61189 448906 61755
rect 1066 60101 448906 60667
rect 1066 59013 448906 59579
rect 1066 57925 448906 58491
rect 1066 56837 448906 57403
rect 1066 55749 448906 56315
rect 1066 54661 448906 55227
rect 1066 53573 448906 54139
rect 1066 52485 448906 53051
rect 1066 51397 448906 51963
rect 1066 50309 448906 50875
rect 1066 49221 448906 49787
rect 1066 48133 448906 48699
rect 1066 47045 448906 47611
rect 1066 45957 448906 46523
rect 1066 44869 448906 45435
rect 1066 43781 448906 44347
rect 1066 42693 448906 43259
rect 1066 41605 448906 42171
rect 1066 40517 448906 41083
rect 1066 39429 448906 39995
rect 1066 38341 448906 38907
rect 1066 37253 448906 37819
rect 1066 36165 448906 36731
rect 1066 35077 448906 35643
rect 1066 33989 448906 34555
rect 1066 32901 448906 33467
rect 1066 31813 448906 32379
rect 1066 30725 448906 31291
rect 1066 29637 448906 30203
rect 1066 28549 448906 29115
rect 1066 27461 448906 28027
rect 1066 26373 448906 26939
rect 1066 25285 448906 25851
rect 1066 24197 448906 24763
rect 1066 23109 448906 23675
rect 1066 22021 448906 22587
rect 1066 20933 448906 21499
rect 1066 19845 448906 20411
rect 1066 18757 448906 19323
rect 1066 17669 448906 18235
rect 1066 16581 448906 17147
rect 1066 15493 448906 16059
rect 1066 14405 448906 14971
rect 1066 13317 448906 13883
rect 1066 12229 448906 12795
rect 1066 11141 448906 11707
rect 1066 10053 448906 10619
rect 1066 8965 448906 9531
rect 1066 7877 448906 8443
rect 1066 6789 448906 7355
rect 1066 5701 448906 6267
rect 1066 4613 448906 5179
rect 1066 3525 448906 4091
rect 1066 2437 448906 3003
<< obsli1 >>
rect 1104 2159 448868 447729
<< obsm1 >>
rect 1104 1980 448868 447760
<< metal2 >>
rect 21270 0 21326 800
rect 22098 0 22154 800
rect 22926 0 22982 800
rect 23754 0 23810 800
rect 24582 0 24638 800
rect 25410 0 25466 800
rect 26238 0 26294 800
rect 27066 0 27122 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30378 0 30434 800
rect 31206 0 31262 800
rect 32034 0 32090 800
rect 32862 0 32918 800
rect 33690 0 33746 800
rect 34518 0 34574 800
rect 35346 0 35402 800
rect 36174 0 36230 800
rect 37002 0 37058 800
rect 37830 0 37886 800
rect 38658 0 38714 800
rect 39486 0 39542 800
rect 40314 0 40370 800
rect 41142 0 41198 800
rect 41970 0 42026 800
rect 42798 0 42854 800
rect 43626 0 43682 800
rect 44454 0 44510 800
rect 45282 0 45338 800
rect 46110 0 46166 800
rect 46938 0 46994 800
rect 47766 0 47822 800
rect 48594 0 48650 800
rect 49422 0 49478 800
rect 50250 0 50306 800
rect 51078 0 51134 800
rect 51906 0 51962 800
rect 52734 0 52790 800
rect 53562 0 53618 800
rect 54390 0 54446 800
rect 55218 0 55274 800
rect 56046 0 56102 800
rect 56874 0 56930 800
rect 57702 0 57758 800
rect 58530 0 58586 800
rect 59358 0 59414 800
rect 60186 0 60242 800
rect 61014 0 61070 800
rect 61842 0 61898 800
rect 62670 0 62726 800
rect 63498 0 63554 800
rect 64326 0 64382 800
rect 65154 0 65210 800
rect 65982 0 66038 800
rect 66810 0 66866 800
rect 67638 0 67694 800
rect 68466 0 68522 800
rect 69294 0 69350 800
rect 70122 0 70178 800
rect 70950 0 71006 800
rect 71778 0 71834 800
rect 72606 0 72662 800
rect 73434 0 73490 800
rect 74262 0 74318 800
rect 75090 0 75146 800
rect 75918 0 75974 800
rect 76746 0 76802 800
rect 77574 0 77630 800
rect 78402 0 78458 800
rect 79230 0 79286 800
rect 80058 0 80114 800
rect 80886 0 80942 800
rect 81714 0 81770 800
rect 82542 0 82598 800
rect 83370 0 83426 800
rect 84198 0 84254 800
rect 85026 0 85082 800
rect 85854 0 85910 800
rect 86682 0 86738 800
rect 87510 0 87566 800
rect 88338 0 88394 800
rect 89166 0 89222 800
rect 89994 0 90050 800
rect 90822 0 90878 800
rect 91650 0 91706 800
rect 92478 0 92534 800
rect 93306 0 93362 800
rect 94134 0 94190 800
rect 94962 0 95018 800
rect 95790 0 95846 800
rect 96618 0 96674 800
rect 97446 0 97502 800
rect 98274 0 98330 800
rect 99102 0 99158 800
rect 99930 0 99986 800
rect 100758 0 100814 800
rect 101586 0 101642 800
rect 102414 0 102470 800
rect 103242 0 103298 800
rect 104070 0 104126 800
rect 104898 0 104954 800
rect 105726 0 105782 800
rect 106554 0 106610 800
rect 107382 0 107438 800
rect 108210 0 108266 800
rect 109038 0 109094 800
rect 109866 0 109922 800
rect 110694 0 110750 800
rect 111522 0 111578 800
rect 112350 0 112406 800
rect 113178 0 113234 800
rect 114006 0 114062 800
rect 114834 0 114890 800
rect 115662 0 115718 800
rect 116490 0 116546 800
rect 117318 0 117374 800
rect 118146 0 118202 800
rect 118974 0 119030 800
rect 119802 0 119858 800
rect 120630 0 120686 800
rect 121458 0 121514 800
rect 122286 0 122342 800
rect 123114 0 123170 800
rect 123942 0 123998 800
rect 124770 0 124826 800
rect 125598 0 125654 800
rect 126426 0 126482 800
rect 127254 0 127310 800
rect 128082 0 128138 800
rect 128910 0 128966 800
rect 129738 0 129794 800
rect 130566 0 130622 800
rect 131394 0 131450 800
rect 132222 0 132278 800
rect 133050 0 133106 800
rect 133878 0 133934 800
rect 134706 0 134762 800
rect 135534 0 135590 800
rect 136362 0 136418 800
rect 137190 0 137246 800
rect 138018 0 138074 800
rect 138846 0 138902 800
rect 139674 0 139730 800
rect 140502 0 140558 800
rect 141330 0 141386 800
rect 142158 0 142214 800
rect 142986 0 143042 800
rect 143814 0 143870 800
rect 144642 0 144698 800
rect 145470 0 145526 800
rect 146298 0 146354 800
rect 147126 0 147182 800
rect 147954 0 148010 800
rect 148782 0 148838 800
rect 149610 0 149666 800
rect 150438 0 150494 800
rect 151266 0 151322 800
rect 152094 0 152150 800
rect 152922 0 152978 800
rect 153750 0 153806 800
rect 154578 0 154634 800
rect 155406 0 155462 800
rect 156234 0 156290 800
rect 157062 0 157118 800
rect 157890 0 157946 800
rect 158718 0 158774 800
rect 159546 0 159602 800
rect 160374 0 160430 800
rect 161202 0 161258 800
rect 162030 0 162086 800
rect 162858 0 162914 800
rect 163686 0 163742 800
rect 164514 0 164570 800
rect 165342 0 165398 800
rect 166170 0 166226 800
rect 166998 0 167054 800
rect 167826 0 167882 800
rect 168654 0 168710 800
rect 169482 0 169538 800
rect 170310 0 170366 800
rect 171138 0 171194 800
rect 171966 0 172022 800
rect 172794 0 172850 800
rect 173622 0 173678 800
rect 174450 0 174506 800
rect 175278 0 175334 800
rect 176106 0 176162 800
rect 176934 0 176990 800
rect 177762 0 177818 800
rect 178590 0 178646 800
rect 179418 0 179474 800
rect 180246 0 180302 800
rect 181074 0 181130 800
rect 181902 0 181958 800
rect 182730 0 182786 800
rect 183558 0 183614 800
rect 184386 0 184442 800
rect 185214 0 185270 800
rect 186042 0 186098 800
rect 186870 0 186926 800
rect 187698 0 187754 800
rect 188526 0 188582 800
rect 189354 0 189410 800
rect 190182 0 190238 800
rect 191010 0 191066 800
rect 191838 0 191894 800
rect 192666 0 192722 800
rect 193494 0 193550 800
rect 194322 0 194378 800
rect 195150 0 195206 800
rect 195978 0 196034 800
rect 196806 0 196862 800
rect 197634 0 197690 800
rect 198462 0 198518 800
rect 199290 0 199346 800
rect 200118 0 200174 800
rect 200946 0 201002 800
rect 201774 0 201830 800
rect 202602 0 202658 800
rect 203430 0 203486 800
rect 204258 0 204314 800
rect 205086 0 205142 800
rect 205914 0 205970 800
rect 206742 0 206798 800
rect 207570 0 207626 800
rect 208398 0 208454 800
rect 209226 0 209282 800
rect 210054 0 210110 800
rect 210882 0 210938 800
rect 211710 0 211766 800
rect 212538 0 212594 800
rect 213366 0 213422 800
rect 214194 0 214250 800
rect 215022 0 215078 800
rect 215850 0 215906 800
rect 216678 0 216734 800
rect 217506 0 217562 800
rect 218334 0 218390 800
rect 219162 0 219218 800
rect 219990 0 220046 800
rect 220818 0 220874 800
rect 221646 0 221702 800
rect 222474 0 222530 800
rect 223302 0 223358 800
rect 224130 0 224186 800
rect 224958 0 225014 800
rect 225786 0 225842 800
rect 226614 0 226670 800
rect 227442 0 227498 800
rect 228270 0 228326 800
rect 229098 0 229154 800
rect 229926 0 229982 800
rect 230754 0 230810 800
rect 231582 0 231638 800
rect 232410 0 232466 800
rect 233238 0 233294 800
rect 234066 0 234122 800
rect 234894 0 234950 800
rect 235722 0 235778 800
rect 236550 0 236606 800
rect 237378 0 237434 800
rect 238206 0 238262 800
rect 239034 0 239090 800
rect 239862 0 239918 800
rect 240690 0 240746 800
rect 241518 0 241574 800
rect 242346 0 242402 800
rect 243174 0 243230 800
rect 244002 0 244058 800
rect 244830 0 244886 800
rect 245658 0 245714 800
rect 246486 0 246542 800
rect 247314 0 247370 800
rect 248142 0 248198 800
rect 248970 0 249026 800
rect 249798 0 249854 800
rect 250626 0 250682 800
rect 251454 0 251510 800
rect 252282 0 252338 800
rect 253110 0 253166 800
rect 253938 0 253994 800
rect 254766 0 254822 800
rect 255594 0 255650 800
rect 256422 0 256478 800
rect 257250 0 257306 800
rect 258078 0 258134 800
rect 258906 0 258962 800
rect 259734 0 259790 800
rect 260562 0 260618 800
rect 261390 0 261446 800
rect 262218 0 262274 800
rect 263046 0 263102 800
rect 263874 0 263930 800
rect 264702 0 264758 800
rect 265530 0 265586 800
rect 266358 0 266414 800
rect 267186 0 267242 800
rect 268014 0 268070 800
rect 268842 0 268898 800
rect 269670 0 269726 800
rect 270498 0 270554 800
rect 271326 0 271382 800
rect 272154 0 272210 800
rect 272982 0 273038 800
rect 273810 0 273866 800
rect 274638 0 274694 800
rect 275466 0 275522 800
rect 276294 0 276350 800
rect 277122 0 277178 800
rect 277950 0 278006 800
rect 278778 0 278834 800
rect 279606 0 279662 800
rect 280434 0 280490 800
rect 281262 0 281318 800
rect 282090 0 282146 800
rect 282918 0 282974 800
rect 283746 0 283802 800
rect 284574 0 284630 800
rect 285402 0 285458 800
rect 286230 0 286286 800
rect 287058 0 287114 800
rect 287886 0 287942 800
rect 288714 0 288770 800
rect 289542 0 289598 800
rect 290370 0 290426 800
rect 291198 0 291254 800
rect 292026 0 292082 800
rect 292854 0 292910 800
rect 293682 0 293738 800
rect 294510 0 294566 800
rect 295338 0 295394 800
rect 296166 0 296222 800
rect 296994 0 297050 800
rect 297822 0 297878 800
rect 298650 0 298706 800
rect 299478 0 299534 800
rect 300306 0 300362 800
rect 301134 0 301190 800
rect 301962 0 302018 800
rect 302790 0 302846 800
rect 303618 0 303674 800
rect 304446 0 304502 800
rect 305274 0 305330 800
rect 306102 0 306158 800
rect 306930 0 306986 800
rect 307758 0 307814 800
rect 308586 0 308642 800
rect 309414 0 309470 800
rect 310242 0 310298 800
rect 311070 0 311126 800
rect 311898 0 311954 800
rect 312726 0 312782 800
rect 313554 0 313610 800
rect 314382 0 314438 800
rect 315210 0 315266 800
rect 316038 0 316094 800
rect 316866 0 316922 800
rect 317694 0 317750 800
rect 318522 0 318578 800
rect 319350 0 319406 800
rect 320178 0 320234 800
rect 321006 0 321062 800
rect 321834 0 321890 800
rect 322662 0 322718 800
rect 323490 0 323546 800
rect 324318 0 324374 800
rect 325146 0 325202 800
rect 325974 0 326030 800
rect 326802 0 326858 800
rect 327630 0 327686 800
rect 328458 0 328514 800
rect 329286 0 329342 800
rect 330114 0 330170 800
rect 330942 0 330998 800
rect 331770 0 331826 800
rect 332598 0 332654 800
rect 333426 0 333482 800
rect 334254 0 334310 800
rect 335082 0 335138 800
rect 335910 0 335966 800
rect 336738 0 336794 800
rect 337566 0 337622 800
rect 338394 0 338450 800
rect 339222 0 339278 800
rect 340050 0 340106 800
rect 340878 0 340934 800
rect 341706 0 341762 800
rect 342534 0 342590 800
rect 343362 0 343418 800
rect 344190 0 344246 800
rect 345018 0 345074 800
rect 345846 0 345902 800
rect 346674 0 346730 800
rect 347502 0 347558 800
rect 348330 0 348386 800
rect 349158 0 349214 800
rect 349986 0 350042 800
rect 350814 0 350870 800
rect 351642 0 351698 800
rect 352470 0 352526 800
rect 353298 0 353354 800
rect 354126 0 354182 800
rect 354954 0 355010 800
rect 355782 0 355838 800
rect 356610 0 356666 800
rect 357438 0 357494 800
rect 358266 0 358322 800
rect 359094 0 359150 800
rect 359922 0 359978 800
rect 360750 0 360806 800
rect 361578 0 361634 800
rect 362406 0 362462 800
rect 363234 0 363290 800
rect 364062 0 364118 800
rect 364890 0 364946 800
rect 365718 0 365774 800
rect 366546 0 366602 800
rect 367374 0 367430 800
rect 368202 0 368258 800
rect 369030 0 369086 800
rect 369858 0 369914 800
rect 370686 0 370742 800
rect 371514 0 371570 800
rect 372342 0 372398 800
rect 373170 0 373226 800
rect 373998 0 374054 800
rect 374826 0 374882 800
rect 375654 0 375710 800
rect 376482 0 376538 800
rect 377310 0 377366 800
rect 378138 0 378194 800
rect 378966 0 379022 800
rect 379794 0 379850 800
rect 380622 0 380678 800
rect 381450 0 381506 800
rect 382278 0 382334 800
rect 383106 0 383162 800
rect 383934 0 383990 800
rect 384762 0 384818 800
rect 385590 0 385646 800
rect 386418 0 386474 800
rect 387246 0 387302 800
rect 388074 0 388130 800
rect 388902 0 388958 800
rect 389730 0 389786 800
rect 390558 0 390614 800
rect 391386 0 391442 800
rect 392214 0 392270 800
rect 393042 0 393098 800
rect 393870 0 393926 800
rect 394698 0 394754 800
rect 395526 0 395582 800
rect 396354 0 396410 800
rect 397182 0 397238 800
rect 398010 0 398066 800
rect 398838 0 398894 800
rect 399666 0 399722 800
rect 400494 0 400550 800
rect 401322 0 401378 800
rect 402150 0 402206 800
rect 402978 0 403034 800
rect 403806 0 403862 800
rect 404634 0 404690 800
rect 405462 0 405518 800
rect 406290 0 406346 800
rect 407118 0 407174 800
rect 407946 0 408002 800
rect 408774 0 408830 800
rect 409602 0 409658 800
rect 410430 0 410486 800
rect 411258 0 411314 800
rect 412086 0 412142 800
rect 412914 0 412970 800
rect 413742 0 413798 800
rect 414570 0 414626 800
rect 415398 0 415454 800
rect 416226 0 416282 800
rect 417054 0 417110 800
rect 417882 0 417938 800
rect 418710 0 418766 800
rect 419538 0 419594 800
rect 420366 0 420422 800
rect 421194 0 421250 800
rect 422022 0 422078 800
rect 422850 0 422906 800
rect 423678 0 423734 800
rect 424506 0 424562 800
rect 425334 0 425390 800
rect 426162 0 426218 800
rect 426990 0 427046 800
rect 427818 0 427874 800
rect 428646 0 428702 800
<< obsm2 >>
rect 1584 856 434602 447749
rect 1584 734 21214 856
rect 21382 734 22042 856
rect 22210 734 22870 856
rect 23038 734 23698 856
rect 23866 734 24526 856
rect 24694 734 25354 856
rect 25522 734 26182 856
rect 26350 734 27010 856
rect 27178 734 27838 856
rect 28006 734 28666 856
rect 28834 734 29494 856
rect 29662 734 30322 856
rect 30490 734 31150 856
rect 31318 734 31978 856
rect 32146 734 32806 856
rect 32974 734 33634 856
rect 33802 734 34462 856
rect 34630 734 35290 856
rect 35458 734 36118 856
rect 36286 734 36946 856
rect 37114 734 37774 856
rect 37942 734 38602 856
rect 38770 734 39430 856
rect 39598 734 40258 856
rect 40426 734 41086 856
rect 41254 734 41914 856
rect 42082 734 42742 856
rect 42910 734 43570 856
rect 43738 734 44398 856
rect 44566 734 45226 856
rect 45394 734 46054 856
rect 46222 734 46882 856
rect 47050 734 47710 856
rect 47878 734 48538 856
rect 48706 734 49366 856
rect 49534 734 50194 856
rect 50362 734 51022 856
rect 51190 734 51850 856
rect 52018 734 52678 856
rect 52846 734 53506 856
rect 53674 734 54334 856
rect 54502 734 55162 856
rect 55330 734 55990 856
rect 56158 734 56818 856
rect 56986 734 57646 856
rect 57814 734 58474 856
rect 58642 734 59302 856
rect 59470 734 60130 856
rect 60298 734 60958 856
rect 61126 734 61786 856
rect 61954 734 62614 856
rect 62782 734 63442 856
rect 63610 734 64270 856
rect 64438 734 65098 856
rect 65266 734 65926 856
rect 66094 734 66754 856
rect 66922 734 67582 856
rect 67750 734 68410 856
rect 68578 734 69238 856
rect 69406 734 70066 856
rect 70234 734 70894 856
rect 71062 734 71722 856
rect 71890 734 72550 856
rect 72718 734 73378 856
rect 73546 734 74206 856
rect 74374 734 75034 856
rect 75202 734 75862 856
rect 76030 734 76690 856
rect 76858 734 77518 856
rect 77686 734 78346 856
rect 78514 734 79174 856
rect 79342 734 80002 856
rect 80170 734 80830 856
rect 80998 734 81658 856
rect 81826 734 82486 856
rect 82654 734 83314 856
rect 83482 734 84142 856
rect 84310 734 84970 856
rect 85138 734 85798 856
rect 85966 734 86626 856
rect 86794 734 87454 856
rect 87622 734 88282 856
rect 88450 734 89110 856
rect 89278 734 89938 856
rect 90106 734 90766 856
rect 90934 734 91594 856
rect 91762 734 92422 856
rect 92590 734 93250 856
rect 93418 734 94078 856
rect 94246 734 94906 856
rect 95074 734 95734 856
rect 95902 734 96562 856
rect 96730 734 97390 856
rect 97558 734 98218 856
rect 98386 734 99046 856
rect 99214 734 99874 856
rect 100042 734 100702 856
rect 100870 734 101530 856
rect 101698 734 102358 856
rect 102526 734 103186 856
rect 103354 734 104014 856
rect 104182 734 104842 856
rect 105010 734 105670 856
rect 105838 734 106498 856
rect 106666 734 107326 856
rect 107494 734 108154 856
rect 108322 734 108982 856
rect 109150 734 109810 856
rect 109978 734 110638 856
rect 110806 734 111466 856
rect 111634 734 112294 856
rect 112462 734 113122 856
rect 113290 734 113950 856
rect 114118 734 114778 856
rect 114946 734 115606 856
rect 115774 734 116434 856
rect 116602 734 117262 856
rect 117430 734 118090 856
rect 118258 734 118918 856
rect 119086 734 119746 856
rect 119914 734 120574 856
rect 120742 734 121402 856
rect 121570 734 122230 856
rect 122398 734 123058 856
rect 123226 734 123886 856
rect 124054 734 124714 856
rect 124882 734 125542 856
rect 125710 734 126370 856
rect 126538 734 127198 856
rect 127366 734 128026 856
rect 128194 734 128854 856
rect 129022 734 129682 856
rect 129850 734 130510 856
rect 130678 734 131338 856
rect 131506 734 132166 856
rect 132334 734 132994 856
rect 133162 734 133822 856
rect 133990 734 134650 856
rect 134818 734 135478 856
rect 135646 734 136306 856
rect 136474 734 137134 856
rect 137302 734 137962 856
rect 138130 734 138790 856
rect 138958 734 139618 856
rect 139786 734 140446 856
rect 140614 734 141274 856
rect 141442 734 142102 856
rect 142270 734 142930 856
rect 143098 734 143758 856
rect 143926 734 144586 856
rect 144754 734 145414 856
rect 145582 734 146242 856
rect 146410 734 147070 856
rect 147238 734 147898 856
rect 148066 734 148726 856
rect 148894 734 149554 856
rect 149722 734 150382 856
rect 150550 734 151210 856
rect 151378 734 152038 856
rect 152206 734 152866 856
rect 153034 734 153694 856
rect 153862 734 154522 856
rect 154690 734 155350 856
rect 155518 734 156178 856
rect 156346 734 157006 856
rect 157174 734 157834 856
rect 158002 734 158662 856
rect 158830 734 159490 856
rect 159658 734 160318 856
rect 160486 734 161146 856
rect 161314 734 161974 856
rect 162142 734 162802 856
rect 162970 734 163630 856
rect 163798 734 164458 856
rect 164626 734 165286 856
rect 165454 734 166114 856
rect 166282 734 166942 856
rect 167110 734 167770 856
rect 167938 734 168598 856
rect 168766 734 169426 856
rect 169594 734 170254 856
rect 170422 734 171082 856
rect 171250 734 171910 856
rect 172078 734 172738 856
rect 172906 734 173566 856
rect 173734 734 174394 856
rect 174562 734 175222 856
rect 175390 734 176050 856
rect 176218 734 176878 856
rect 177046 734 177706 856
rect 177874 734 178534 856
rect 178702 734 179362 856
rect 179530 734 180190 856
rect 180358 734 181018 856
rect 181186 734 181846 856
rect 182014 734 182674 856
rect 182842 734 183502 856
rect 183670 734 184330 856
rect 184498 734 185158 856
rect 185326 734 185986 856
rect 186154 734 186814 856
rect 186982 734 187642 856
rect 187810 734 188470 856
rect 188638 734 189298 856
rect 189466 734 190126 856
rect 190294 734 190954 856
rect 191122 734 191782 856
rect 191950 734 192610 856
rect 192778 734 193438 856
rect 193606 734 194266 856
rect 194434 734 195094 856
rect 195262 734 195922 856
rect 196090 734 196750 856
rect 196918 734 197578 856
rect 197746 734 198406 856
rect 198574 734 199234 856
rect 199402 734 200062 856
rect 200230 734 200890 856
rect 201058 734 201718 856
rect 201886 734 202546 856
rect 202714 734 203374 856
rect 203542 734 204202 856
rect 204370 734 205030 856
rect 205198 734 205858 856
rect 206026 734 206686 856
rect 206854 734 207514 856
rect 207682 734 208342 856
rect 208510 734 209170 856
rect 209338 734 209998 856
rect 210166 734 210826 856
rect 210994 734 211654 856
rect 211822 734 212482 856
rect 212650 734 213310 856
rect 213478 734 214138 856
rect 214306 734 214966 856
rect 215134 734 215794 856
rect 215962 734 216622 856
rect 216790 734 217450 856
rect 217618 734 218278 856
rect 218446 734 219106 856
rect 219274 734 219934 856
rect 220102 734 220762 856
rect 220930 734 221590 856
rect 221758 734 222418 856
rect 222586 734 223246 856
rect 223414 734 224074 856
rect 224242 734 224902 856
rect 225070 734 225730 856
rect 225898 734 226558 856
rect 226726 734 227386 856
rect 227554 734 228214 856
rect 228382 734 229042 856
rect 229210 734 229870 856
rect 230038 734 230698 856
rect 230866 734 231526 856
rect 231694 734 232354 856
rect 232522 734 233182 856
rect 233350 734 234010 856
rect 234178 734 234838 856
rect 235006 734 235666 856
rect 235834 734 236494 856
rect 236662 734 237322 856
rect 237490 734 238150 856
rect 238318 734 238978 856
rect 239146 734 239806 856
rect 239974 734 240634 856
rect 240802 734 241462 856
rect 241630 734 242290 856
rect 242458 734 243118 856
rect 243286 734 243946 856
rect 244114 734 244774 856
rect 244942 734 245602 856
rect 245770 734 246430 856
rect 246598 734 247258 856
rect 247426 734 248086 856
rect 248254 734 248914 856
rect 249082 734 249742 856
rect 249910 734 250570 856
rect 250738 734 251398 856
rect 251566 734 252226 856
rect 252394 734 253054 856
rect 253222 734 253882 856
rect 254050 734 254710 856
rect 254878 734 255538 856
rect 255706 734 256366 856
rect 256534 734 257194 856
rect 257362 734 258022 856
rect 258190 734 258850 856
rect 259018 734 259678 856
rect 259846 734 260506 856
rect 260674 734 261334 856
rect 261502 734 262162 856
rect 262330 734 262990 856
rect 263158 734 263818 856
rect 263986 734 264646 856
rect 264814 734 265474 856
rect 265642 734 266302 856
rect 266470 734 267130 856
rect 267298 734 267958 856
rect 268126 734 268786 856
rect 268954 734 269614 856
rect 269782 734 270442 856
rect 270610 734 271270 856
rect 271438 734 272098 856
rect 272266 734 272926 856
rect 273094 734 273754 856
rect 273922 734 274582 856
rect 274750 734 275410 856
rect 275578 734 276238 856
rect 276406 734 277066 856
rect 277234 734 277894 856
rect 278062 734 278722 856
rect 278890 734 279550 856
rect 279718 734 280378 856
rect 280546 734 281206 856
rect 281374 734 282034 856
rect 282202 734 282862 856
rect 283030 734 283690 856
rect 283858 734 284518 856
rect 284686 734 285346 856
rect 285514 734 286174 856
rect 286342 734 287002 856
rect 287170 734 287830 856
rect 287998 734 288658 856
rect 288826 734 289486 856
rect 289654 734 290314 856
rect 290482 734 291142 856
rect 291310 734 291970 856
rect 292138 734 292798 856
rect 292966 734 293626 856
rect 293794 734 294454 856
rect 294622 734 295282 856
rect 295450 734 296110 856
rect 296278 734 296938 856
rect 297106 734 297766 856
rect 297934 734 298594 856
rect 298762 734 299422 856
rect 299590 734 300250 856
rect 300418 734 301078 856
rect 301246 734 301906 856
rect 302074 734 302734 856
rect 302902 734 303562 856
rect 303730 734 304390 856
rect 304558 734 305218 856
rect 305386 734 306046 856
rect 306214 734 306874 856
rect 307042 734 307702 856
rect 307870 734 308530 856
rect 308698 734 309358 856
rect 309526 734 310186 856
rect 310354 734 311014 856
rect 311182 734 311842 856
rect 312010 734 312670 856
rect 312838 734 313498 856
rect 313666 734 314326 856
rect 314494 734 315154 856
rect 315322 734 315982 856
rect 316150 734 316810 856
rect 316978 734 317638 856
rect 317806 734 318466 856
rect 318634 734 319294 856
rect 319462 734 320122 856
rect 320290 734 320950 856
rect 321118 734 321778 856
rect 321946 734 322606 856
rect 322774 734 323434 856
rect 323602 734 324262 856
rect 324430 734 325090 856
rect 325258 734 325918 856
rect 326086 734 326746 856
rect 326914 734 327574 856
rect 327742 734 328402 856
rect 328570 734 329230 856
rect 329398 734 330058 856
rect 330226 734 330886 856
rect 331054 734 331714 856
rect 331882 734 332542 856
rect 332710 734 333370 856
rect 333538 734 334198 856
rect 334366 734 335026 856
rect 335194 734 335854 856
rect 336022 734 336682 856
rect 336850 734 337510 856
rect 337678 734 338338 856
rect 338506 734 339166 856
rect 339334 734 339994 856
rect 340162 734 340822 856
rect 340990 734 341650 856
rect 341818 734 342478 856
rect 342646 734 343306 856
rect 343474 734 344134 856
rect 344302 734 344962 856
rect 345130 734 345790 856
rect 345958 734 346618 856
rect 346786 734 347446 856
rect 347614 734 348274 856
rect 348442 734 349102 856
rect 349270 734 349930 856
rect 350098 734 350758 856
rect 350926 734 351586 856
rect 351754 734 352414 856
rect 352582 734 353242 856
rect 353410 734 354070 856
rect 354238 734 354898 856
rect 355066 734 355726 856
rect 355894 734 356554 856
rect 356722 734 357382 856
rect 357550 734 358210 856
rect 358378 734 359038 856
rect 359206 734 359866 856
rect 360034 734 360694 856
rect 360862 734 361522 856
rect 361690 734 362350 856
rect 362518 734 363178 856
rect 363346 734 364006 856
rect 364174 734 364834 856
rect 365002 734 365662 856
rect 365830 734 366490 856
rect 366658 734 367318 856
rect 367486 734 368146 856
rect 368314 734 368974 856
rect 369142 734 369802 856
rect 369970 734 370630 856
rect 370798 734 371458 856
rect 371626 734 372286 856
rect 372454 734 373114 856
rect 373282 734 373942 856
rect 374110 734 374770 856
rect 374938 734 375598 856
rect 375766 734 376426 856
rect 376594 734 377254 856
rect 377422 734 378082 856
rect 378250 734 378910 856
rect 379078 734 379738 856
rect 379906 734 380566 856
rect 380734 734 381394 856
rect 381562 734 382222 856
rect 382390 734 383050 856
rect 383218 734 383878 856
rect 384046 734 384706 856
rect 384874 734 385534 856
rect 385702 734 386362 856
rect 386530 734 387190 856
rect 387358 734 388018 856
rect 388186 734 388846 856
rect 389014 734 389674 856
rect 389842 734 390502 856
rect 390670 734 391330 856
rect 391498 734 392158 856
rect 392326 734 392986 856
rect 393154 734 393814 856
rect 393982 734 394642 856
rect 394810 734 395470 856
rect 395638 734 396298 856
rect 396466 734 397126 856
rect 397294 734 397954 856
rect 398122 734 398782 856
rect 398950 734 399610 856
rect 399778 734 400438 856
rect 400606 734 401266 856
rect 401434 734 402094 856
rect 402262 734 402922 856
rect 403090 734 403750 856
rect 403918 734 404578 856
rect 404746 734 405406 856
rect 405574 734 406234 856
rect 406402 734 407062 856
rect 407230 734 407890 856
rect 408058 734 408718 856
rect 408886 734 409546 856
rect 409714 734 410374 856
rect 410542 734 411202 856
rect 411370 734 412030 856
rect 412198 734 412858 856
rect 413026 734 413686 856
rect 413854 734 414514 856
rect 414682 734 415342 856
rect 415510 734 416170 856
rect 416338 734 416998 856
rect 417166 734 417826 856
rect 417994 734 418654 856
rect 418822 734 419482 856
rect 419650 734 420310 856
rect 420478 734 421138 856
rect 421306 734 421966 856
rect 422134 734 422794 856
rect 422962 734 423622 856
rect 423790 734 424450 856
rect 424618 734 425278 856
rect 425446 734 426106 856
rect 426274 734 426934 856
rect 427102 734 427762 856
rect 427930 734 428590 856
rect 428758 734 434602 856
<< obsm3 >>
rect 4210 2143 434606 447745
<< metal4 >>
rect 4208 2128 4528 447760
rect 19568 2128 19888 447760
rect 34928 2128 35248 447760
rect 50288 2128 50608 447760
rect 65648 2128 65968 447760
rect 81008 2128 81328 447760
rect 96368 2128 96688 447760
rect 111728 2128 112048 447760
rect 127088 2128 127408 447760
rect 142448 2128 142768 447760
rect 157808 2128 158128 447760
rect 173168 2128 173488 447760
rect 188528 2128 188848 447760
rect 203888 2128 204208 447760
rect 219248 2128 219568 447760
rect 234608 2128 234928 447760
rect 249968 2128 250288 447760
rect 265328 2128 265648 447760
rect 280688 2128 281008 447760
rect 296048 2128 296368 447760
rect 311408 2128 311728 447760
rect 326768 2128 327088 447760
rect 342128 2128 342448 447760
rect 357488 2128 357808 447760
rect 372848 2128 373168 447760
rect 388208 2128 388528 447760
rect 403568 2128 403888 447760
rect 418928 2128 419248 447760
rect 434288 2128 434608 447760
<< obsm4 >>
rect 34651 3299 34848 67285
rect 35328 3299 50208 67285
rect 50688 3299 65568 67285
rect 66048 3299 80928 67285
rect 81408 3299 85685 67285
<< labels >>
rlabel metal2 s 426990 0 427046 800 6 irq[0]
port 1 nsew signal output
rlabel metal2 s 427818 0 427874 800 6 irq[1]
port 2 nsew signal output
rlabel metal2 s 428646 0 428702 800 6 irq[2]
port 3 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_in[0]
port 4 nsew signal input
rlabel metal2 s 357438 0 357494 800 6 la_data_in[100]
port 5 nsew signal input
rlabel metal2 s 359922 0 359978 800 6 la_data_in[101]
port 6 nsew signal input
rlabel metal2 s 362406 0 362462 800 6 la_data_in[102]
port 7 nsew signal input
rlabel metal2 s 364890 0 364946 800 6 la_data_in[103]
port 8 nsew signal input
rlabel metal2 s 367374 0 367430 800 6 la_data_in[104]
port 9 nsew signal input
rlabel metal2 s 369858 0 369914 800 6 la_data_in[105]
port 10 nsew signal input
rlabel metal2 s 372342 0 372398 800 6 la_data_in[106]
port 11 nsew signal input
rlabel metal2 s 374826 0 374882 800 6 la_data_in[107]
port 12 nsew signal input
rlabel metal2 s 377310 0 377366 800 6 la_data_in[108]
port 13 nsew signal input
rlabel metal2 s 379794 0 379850 800 6 la_data_in[109]
port 14 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_data_in[10]
port 15 nsew signal input
rlabel metal2 s 382278 0 382334 800 6 la_data_in[110]
port 16 nsew signal input
rlabel metal2 s 384762 0 384818 800 6 la_data_in[111]
port 17 nsew signal input
rlabel metal2 s 387246 0 387302 800 6 la_data_in[112]
port 18 nsew signal input
rlabel metal2 s 389730 0 389786 800 6 la_data_in[113]
port 19 nsew signal input
rlabel metal2 s 392214 0 392270 800 6 la_data_in[114]
port 20 nsew signal input
rlabel metal2 s 394698 0 394754 800 6 la_data_in[115]
port 21 nsew signal input
rlabel metal2 s 397182 0 397238 800 6 la_data_in[116]
port 22 nsew signal input
rlabel metal2 s 399666 0 399722 800 6 la_data_in[117]
port 23 nsew signal input
rlabel metal2 s 402150 0 402206 800 6 la_data_in[118]
port 24 nsew signal input
rlabel metal2 s 404634 0 404690 800 6 la_data_in[119]
port 25 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_data_in[11]
port 26 nsew signal input
rlabel metal2 s 407118 0 407174 800 6 la_data_in[120]
port 27 nsew signal input
rlabel metal2 s 409602 0 409658 800 6 la_data_in[121]
port 28 nsew signal input
rlabel metal2 s 412086 0 412142 800 6 la_data_in[122]
port 29 nsew signal input
rlabel metal2 s 414570 0 414626 800 6 la_data_in[123]
port 30 nsew signal input
rlabel metal2 s 417054 0 417110 800 6 la_data_in[124]
port 31 nsew signal input
rlabel metal2 s 419538 0 419594 800 6 la_data_in[125]
port 32 nsew signal input
rlabel metal2 s 422022 0 422078 800 6 la_data_in[126]
port 33 nsew signal input
rlabel metal2 s 424506 0 424562 800 6 la_data_in[127]
port 34 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 la_data_in[12]
port 35 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_data_in[13]
port 36 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_data_in[14]
port 37 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 la_data_in[15]
port 38 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_data_in[16]
port 39 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_data_in[17]
port 40 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_data_in[18]
port 41 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_data_in[19]
port 42 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[1]
port 43 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_data_in[20]
port 44 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 la_data_in[21]
port 45 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 la_data_in[22]
port 46 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_data_in[23]
port 47 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_data_in[24]
port 48 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 la_data_in[25]
port 49 nsew signal input
rlabel metal2 s 173622 0 173678 800 6 la_data_in[26]
port 50 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_data_in[27]
port 51 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_data_in[28]
port 52 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 la_data_in[29]
port 53 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[2]
port 54 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 la_data_in[30]
port 55 nsew signal input
rlabel metal2 s 186042 0 186098 800 6 la_data_in[31]
port 56 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_data_in[32]
port 57 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 la_data_in[33]
port 58 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_data_in[34]
port 59 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 la_data_in[35]
port 60 nsew signal input
rlabel metal2 s 198462 0 198518 800 6 la_data_in[36]
port 61 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 la_data_in[37]
port 62 nsew signal input
rlabel metal2 s 203430 0 203486 800 6 la_data_in[38]
port 63 nsew signal input
rlabel metal2 s 205914 0 205970 800 6 la_data_in[39]
port 64 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_data_in[3]
port 65 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_data_in[40]
port 66 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_data_in[41]
port 67 nsew signal input
rlabel metal2 s 213366 0 213422 800 6 la_data_in[42]
port 68 nsew signal input
rlabel metal2 s 215850 0 215906 800 6 la_data_in[43]
port 69 nsew signal input
rlabel metal2 s 218334 0 218390 800 6 la_data_in[44]
port 70 nsew signal input
rlabel metal2 s 220818 0 220874 800 6 la_data_in[45]
port 71 nsew signal input
rlabel metal2 s 223302 0 223358 800 6 la_data_in[46]
port 72 nsew signal input
rlabel metal2 s 225786 0 225842 800 6 la_data_in[47]
port 73 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_data_in[48]
port 74 nsew signal input
rlabel metal2 s 230754 0 230810 800 6 la_data_in[49]
port 75 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[4]
port 76 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_data_in[50]
port 77 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_data_in[51]
port 78 nsew signal input
rlabel metal2 s 238206 0 238262 800 6 la_data_in[52]
port 79 nsew signal input
rlabel metal2 s 240690 0 240746 800 6 la_data_in[53]
port 80 nsew signal input
rlabel metal2 s 243174 0 243230 800 6 la_data_in[54]
port 81 nsew signal input
rlabel metal2 s 245658 0 245714 800 6 la_data_in[55]
port 82 nsew signal input
rlabel metal2 s 248142 0 248198 800 6 la_data_in[56]
port 83 nsew signal input
rlabel metal2 s 250626 0 250682 800 6 la_data_in[57]
port 84 nsew signal input
rlabel metal2 s 253110 0 253166 800 6 la_data_in[58]
port 85 nsew signal input
rlabel metal2 s 255594 0 255650 800 6 la_data_in[59]
port 86 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 la_data_in[5]
port 87 nsew signal input
rlabel metal2 s 258078 0 258134 800 6 la_data_in[60]
port 88 nsew signal input
rlabel metal2 s 260562 0 260618 800 6 la_data_in[61]
port 89 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_data_in[62]
port 90 nsew signal input
rlabel metal2 s 265530 0 265586 800 6 la_data_in[63]
port 91 nsew signal input
rlabel metal2 s 268014 0 268070 800 6 la_data_in[64]
port 92 nsew signal input
rlabel metal2 s 270498 0 270554 800 6 la_data_in[65]
port 93 nsew signal input
rlabel metal2 s 272982 0 273038 800 6 la_data_in[66]
port 94 nsew signal input
rlabel metal2 s 275466 0 275522 800 6 la_data_in[67]
port 95 nsew signal input
rlabel metal2 s 277950 0 278006 800 6 la_data_in[68]
port 96 nsew signal input
rlabel metal2 s 280434 0 280490 800 6 la_data_in[69]
port 97 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_data_in[6]
port 98 nsew signal input
rlabel metal2 s 282918 0 282974 800 6 la_data_in[70]
port 99 nsew signal input
rlabel metal2 s 285402 0 285458 800 6 la_data_in[71]
port 100 nsew signal input
rlabel metal2 s 287886 0 287942 800 6 la_data_in[72]
port 101 nsew signal input
rlabel metal2 s 290370 0 290426 800 6 la_data_in[73]
port 102 nsew signal input
rlabel metal2 s 292854 0 292910 800 6 la_data_in[74]
port 103 nsew signal input
rlabel metal2 s 295338 0 295394 800 6 la_data_in[75]
port 104 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_data_in[76]
port 105 nsew signal input
rlabel metal2 s 300306 0 300362 800 6 la_data_in[77]
port 106 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_data_in[78]
port 107 nsew signal input
rlabel metal2 s 305274 0 305330 800 6 la_data_in[79]
port 108 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[7]
port 109 nsew signal input
rlabel metal2 s 307758 0 307814 800 6 la_data_in[80]
port 110 nsew signal input
rlabel metal2 s 310242 0 310298 800 6 la_data_in[81]
port 111 nsew signal input
rlabel metal2 s 312726 0 312782 800 6 la_data_in[82]
port 112 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_data_in[83]
port 113 nsew signal input
rlabel metal2 s 317694 0 317750 800 6 la_data_in[84]
port 114 nsew signal input
rlabel metal2 s 320178 0 320234 800 6 la_data_in[85]
port 115 nsew signal input
rlabel metal2 s 322662 0 322718 800 6 la_data_in[86]
port 116 nsew signal input
rlabel metal2 s 325146 0 325202 800 6 la_data_in[87]
port 117 nsew signal input
rlabel metal2 s 327630 0 327686 800 6 la_data_in[88]
port 118 nsew signal input
rlabel metal2 s 330114 0 330170 800 6 la_data_in[89]
port 119 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[8]
port 120 nsew signal input
rlabel metal2 s 332598 0 332654 800 6 la_data_in[90]
port 121 nsew signal input
rlabel metal2 s 335082 0 335138 800 6 la_data_in[91]
port 122 nsew signal input
rlabel metal2 s 337566 0 337622 800 6 la_data_in[92]
port 123 nsew signal input
rlabel metal2 s 340050 0 340106 800 6 la_data_in[93]
port 124 nsew signal input
rlabel metal2 s 342534 0 342590 800 6 la_data_in[94]
port 125 nsew signal input
rlabel metal2 s 345018 0 345074 800 6 la_data_in[95]
port 126 nsew signal input
rlabel metal2 s 347502 0 347558 800 6 la_data_in[96]
port 127 nsew signal input
rlabel metal2 s 349986 0 350042 800 6 la_data_in[97]
port 128 nsew signal input
rlabel metal2 s 352470 0 352526 800 6 la_data_in[98]
port 129 nsew signal input
rlabel metal2 s 354954 0 355010 800 6 la_data_in[99]
port 130 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[9]
port 131 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_data_out[0]
port 132 nsew signal output
rlabel metal2 s 358266 0 358322 800 6 la_data_out[100]
port 133 nsew signal output
rlabel metal2 s 360750 0 360806 800 6 la_data_out[101]
port 134 nsew signal output
rlabel metal2 s 363234 0 363290 800 6 la_data_out[102]
port 135 nsew signal output
rlabel metal2 s 365718 0 365774 800 6 la_data_out[103]
port 136 nsew signal output
rlabel metal2 s 368202 0 368258 800 6 la_data_out[104]
port 137 nsew signal output
rlabel metal2 s 370686 0 370742 800 6 la_data_out[105]
port 138 nsew signal output
rlabel metal2 s 373170 0 373226 800 6 la_data_out[106]
port 139 nsew signal output
rlabel metal2 s 375654 0 375710 800 6 la_data_out[107]
port 140 nsew signal output
rlabel metal2 s 378138 0 378194 800 6 la_data_out[108]
port 141 nsew signal output
rlabel metal2 s 380622 0 380678 800 6 la_data_out[109]
port 142 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 la_data_out[10]
port 143 nsew signal output
rlabel metal2 s 383106 0 383162 800 6 la_data_out[110]
port 144 nsew signal output
rlabel metal2 s 385590 0 385646 800 6 la_data_out[111]
port 145 nsew signal output
rlabel metal2 s 388074 0 388130 800 6 la_data_out[112]
port 146 nsew signal output
rlabel metal2 s 390558 0 390614 800 6 la_data_out[113]
port 147 nsew signal output
rlabel metal2 s 393042 0 393098 800 6 la_data_out[114]
port 148 nsew signal output
rlabel metal2 s 395526 0 395582 800 6 la_data_out[115]
port 149 nsew signal output
rlabel metal2 s 398010 0 398066 800 6 la_data_out[116]
port 150 nsew signal output
rlabel metal2 s 400494 0 400550 800 6 la_data_out[117]
port 151 nsew signal output
rlabel metal2 s 402978 0 403034 800 6 la_data_out[118]
port 152 nsew signal output
rlabel metal2 s 405462 0 405518 800 6 la_data_out[119]
port 153 nsew signal output
rlabel metal2 s 137190 0 137246 800 6 la_data_out[11]
port 154 nsew signal output
rlabel metal2 s 407946 0 408002 800 6 la_data_out[120]
port 155 nsew signal output
rlabel metal2 s 410430 0 410486 800 6 la_data_out[121]
port 156 nsew signal output
rlabel metal2 s 412914 0 412970 800 6 la_data_out[122]
port 157 nsew signal output
rlabel metal2 s 415398 0 415454 800 6 la_data_out[123]
port 158 nsew signal output
rlabel metal2 s 417882 0 417938 800 6 la_data_out[124]
port 159 nsew signal output
rlabel metal2 s 420366 0 420422 800 6 la_data_out[125]
port 160 nsew signal output
rlabel metal2 s 422850 0 422906 800 6 la_data_out[126]
port 161 nsew signal output
rlabel metal2 s 425334 0 425390 800 6 la_data_out[127]
port 162 nsew signal output
rlabel metal2 s 139674 0 139730 800 6 la_data_out[12]
port 163 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 la_data_out[13]
port 164 nsew signal output
rlabel metal2 s 144642 0 144698 800 6 la_data_out[14]
port 165 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 la_data_out[15]
port 166 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[16]
port 167 nsew signal output
rlabel metal2 s 152094 0 152150 800 6 la_data_out[17]
port 168 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 la_data_out[18]
port 169 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[19]
port 170 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 la_data_out[1]
port 171 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[20]
port 172 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 la_data_out[21]
port 173 nsew signal output
rlabel metal2 s 164514 0 164570 800 6 la_data_out[22]
port 174 nsew signal output
rlabel metal2 s 166998 0 167054 800 6 la_data_out[23]
port 175 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[24]
port 176 nsew signal output
rlabel metal2 s 171966 0 172022 800 6 la_data_out[25]
port 177 nsew signal output
rlabel metal2 s 174450 0 174506 800 6 la_data_out[26]
port 178 nsew signal output
rlabel metal2 s 176934 0 176990 800 6 la_data_out[27]
port 179 nsew signal output
rlabel metal2 s 179418 0 179474 800 6 la_data_out[28]
port 180 nsew signal output
rlabel metal2 s 181902 0 181958 800 6 la_data_out[29]
port 181 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[2]
port 182 nsew signal output
rlabel metal2 s 184386 0 184442 800 6 la_data_out[30]
port 183 nsew signal output
rlabel metal2 s 186870 0 186926 800 6 la_data_out[31]
port 184 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 la_data_out[32]
port 185 nsew signal output
rlabel metal2 s 191838 0 191894 800 6 la_data_out[33]
port 186 nsew signal output
rlabel metal2 s 194322 0 194378 800 6 la_data_out[34]
port 187 nsew signal output
rlabel metal2 s 196806 0 196862 800 6 la_data_out[35]
port 188 nsew signal output
rlabel metal2 s 199290 0 199346 800 6 la_data_out[36]
port 189 nsew signal output
rlabel metal2 s 201774 0 201830 800 6 la_data_out[37]
port 190 nsew signal output
rlabel metal2 s 204258 0 204314 800 6 la_data_out[38]
port 191 nsew signal output
rlabel metal2 s 206742 0 206798 800 6 la_data_out[39]
port 192 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 la_data_out[3]
port 193 nsew signal output
rlabel metal2 s 209226 0 209282 800 6 la_data_out[40]
port 194 nsew signal output
rlabel metal2 s 211710 0 211766 800 6 la_data_out[41]
port 195 nsew signal output
rlabel metal2 s 214194 0 214250 800 6 la_data_out[42]
port 196 nsew signal output
rlabel metal2 s 216678 0 216734 800 6 la_data_out[43]
port 197 nsew signal output
rlabel metal2 s 219162 0 219218 800 6 la_data_out[44]
port 198 nsew signal output
rlabel metal2 s 221646 0 221702 800 6 la_data_out[45]
port 199 nsew signal output
rlabel metal2 s 224130 0 224186 800 6 la_data_out[46]
port 200 nsew signal output
rlabel metal2 s 226614 0 226670 800 6 la_data_out[47]
port 201 nsew signal output
rlabel metal2 s 229098 0 229154 800 6 la_data_out[48]
port 202 nsew signal output
rlabel metal2 s 231582 0 231638 800 6 la_data_out[49]
port 203 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 la_data_out[4]
port 204 nsew signal output
rlabel metal2 s 234066 0 234122 800 6 la_data_out[50]
port 205 nsew signal output
rlabel metal2 s 236550 0 236606 800 6 la_data_out[51]
port 206 nsew signal output
rlabel metal2 s 239034 0 239090 800 6 la_data_out[52]
port 207 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 la_data_out[53]
port 208 nsew signal output
rlabel metal2 s 244002 0 244058 800 6 la_data_out[54]
port 209 nsew signal output
rlabel metal2 s 246486 0 246542 800 6 la_data_out[55]
port 210 nsew signal output
rlabel metal2 s 248970 0 249026 800 6 la_data_out[56]
port 211 nsew signal output
rlabel metal2 s 251454 0 251510 800 6 la_data_out[57]
port 212 nsew signal output
rlabel metal2 s 253938 0 253994 800 6 la_data_out[58]
port 213 nsew signal output
rlabel metal2 s 256422 0 256478 800 6 la_data_out[59]
port 214 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[5]
port 215 nsew signal output
rlabel metal2 s 258906 0 258962 800 6 la_data_out[60]
port 216 nsew signal output
rlabel metal2 s 261390 0 261446 800 6 la_data_out[61]
port 217 nsew signal output
rlabel metal2 s 263874 0 263930 800 6 la_data_out[62]
port 218 nsew signal output
rlabel metal2 s 266358 0 266414 800 6 la_data_out[63]
port 219 nsew signal output
rlabel metal2 s 268842 0 268898 800 6 la_data_out[64]
port 220 nsew signal output
rlabel metal2 s 271326 0 271382 800 6 la_data_out[65]
port 221 nsew signal output
rlabel metal2 s 273810 0 273866 800 6 la_data_out[66]
port 222 nsew signal output
rlabel metal2 s 276294 0 276350 800 6 la_data_out[67]
port 223 nsew signal output
rlabel metal2 s 278778 0 278834 800 6 la_data_out[68]
port 224 nsew signal output
rlabel metal2 s 281262 0 281318 800 6 la_data_out[69]
port 225 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 la_data_out[6]
port 226 nsew signal output
rlabel metal2 s 283746 0 283802 800 6 la_data_out[70]
port 227 nsew signal output
rlabel metal2 s 286230 0 286286 800 6 la_data_out[71]
port 228 nsew signal output
rlabel metal2 s 288714 0 288770 800 6 la_data_out[72]
port 229 nsew signal output
rlabel metal2 s 291198 0 291254 800 6 la_data_out[73]
port 230 nsew signal output
rlabel metal2 s 293682 0 293738 800 6 la_data_out[74]
port 231 nsew signal output
rlabel metal2 s 296166 0 296222 800 6 la_data_out[75]
port 232 nsew signal output
rlabel metal2 s 298650 0 298706 800 6 la_data_out[76]
port 233 nsew signal output
rlabel metal2 s 301134 0 301190 800 6 la_data_out[77]
port 234 nsew signal output
rlabel metal2 s 303618 0 303674 800 6 la_data_out[78]
port 235 nsew signal output
rlabel metal2 s 306102 0 306158 800 6 la_data_out[79]
port 236 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[7]
port 237 nsew signal output
rlabel metal2 s 308586 0 308642 800 6 la_data_out[80]
port 238 nsew signal output
rlabel metal2 s 311070 0 311126 800 6 la_data_out[81]
port 239 nsew signal output
rlabel metal2 s 313554 0 313610 800 6 la_data_out[82]
port 240 nsew signal output
rlabel metal2 s 316038 0 316094 800 6 la_data_out[83]
port 241 nsew signal output
rlabel metal2 s 318522 0 318578 800 6 la_data_out[84]
port 242 nsew signal output
rlabel metal2 s 321006 0 321062 800 6 la_data_out[85]
port 243 nsew signal output
rlabel metal2 s 323490 0 323546 800 6 la_data_out[86]
port 244 nsew signal output
rlabel metal2 s 325974 0 326030 800 6 la_data_out[87]
port 245 nsew signal output
rlabel metal2 s 328458 0 328514 800 6 la_data_out[88]
port 246 nsew signal output
rlabel metal2 s 330942 0 330998 800 6 la_data_out[89]
port 247 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[8]
port 248 nsew signal output
rlabel metal2 s 333426 0 333482 800 6 la_data_out[90]
port 249 nsew signal output
rlabel metal2 s 335910 0 335966 800 6 la_data_out[91]
port 250 nsew signal output
rlabel metal2 s 338394 0 338450 800 6 la_data_out[92]
port 251 nsew signal output
rlabel metal2 s 340878 0 340934 800 6 la_data_out[93]
port 252 nsew signal output
rlabel metal2 s 343362 0 343418 800 6 la_data_out[94]
port 253 nsew signal output
rlabel metal2 s 345846 0 345902 800 6 la_data_out[95]
port 254 nsew signal output
rlabel metal2 s 348330 0 348386 800 6 la_data_out[96]
port 255 nsew signal output
rlabel metal2 s 350814 0 350870 800 6 la_data_out[97]
port 256 nsew signal output
rlabel metal2 s 353298 0 353354 800 6 la_data_out[98]
port 257 nsew signal output
rlabel metal2 s 355782 0 355838 800 6 la_data_out[99]
port 258 nsew signal output
rlabel metal2 s 132222 0 132278 800 6 la_data_out[9]
port 259 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_oenb[0]
port 260 nsew signal input
rlabel metal2 s 359094 0 359150 800 6 la_oenb[100]
port 261 nsew signal input
rlabel metal2 s 361578 0 361634 800 6 la_oenb[101]
port 262 nsew signal input
rlabel metal2 s 364062 0 364118 800 6 la_oenb[102]
port 263 nsew signal input
rlabel metal2 s 366546 0 366602 800 6 la_oenb[103]
port 264 nsew signal input
rlabel metal2 s 369030 0 369086 800 6 la_oenb[104]
port 265 nsew signal input
rlabel metal2 s 371514 0 371570 800 6 la_oenb[105]
port 266 nsew signal input
rlabel metal2 s 373998 0 374054 800 6 la_oenb[106]
port 267 nsew signal input
rlabel metal2 s 376482 0 376538 800 6 la_oenb[107]
port 268 nsew signal input
rlabel metal2 s 378966 0 379022 800 6 la_oenb[108]
port 269 nsew signal input
rlabel metal2 s 381450 0 381506 800 6 la_oenb[109]
port 270 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oenb[10]
port 271 nsew signal input
rlabel metal2 s 383934 0 383990 800 6 la_oenb[110]
port 272 nsew signal input
rlabel metal2 s 386418 0 386474 800 6 la_oenb[111]
port 273 nsew signal input
rlabel metal2 s 388902 0 388958 800 6 la_oenb[112]
port 274 nsew signal input
rlabel metal2 s 391386 0 391442 800 6 la_oenb[113]
port 275 nsew signal input
rlabel metal2 s 393870 0 393926 800 6 la_oenb[114]
port 276 nsew signal input
rlabel metal2 s 396354 0 396410 800 6 la_oenb[115]
port 277 nsew signal input
rlabel metal2 s 398838 0 398894 800 6 la_oenb[116]
port 278 nsew signal input
rlabel metal2 s 401322 0 401378 800 6 la_oenb[117]
port 279 nsew signal input
rlabel metal2 s 403806 0 403862 800 6 la_oenb[118]
port 280 nsew signal input
rlabel metal2 s 406290 0 406346 800 6 la_oenb[119]
port 281 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_oenb[11]
port 282 nsew signal input
rlabel metal2 s 408774 0 408830 800 6 la_oenb[120]
port 283 nsew signal input
rlabel metal2 s 411258 0 411314 800 6 la_oenb[121]
port 284 nsew signal input
rlabel metal2 s 413742 0 413798 800 6 la_oenb[122]
port 285 nsew signal input
rlabel metal2 s 416226 0 416282 800 6 la_oenb[123]
port 286 nsew signal input
rlabel metal2 s 418710 0 418766 800 6 la_oenb[124]
port 287 nsew signal input
rlabel metal2 s 421194 0 421250 800 6 la_oenb[125]
port 288 nsew signal input
rlabel metal2 s 423678 0 423734 800 6 la_oenb[126]
port 289 nsew signal input
rlabel metal2 s 426162 0 426218 800 6 la_oenb[127]
port 290 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 la_oenb[12]
port 291 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_oenb[13]
port 292 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 la_oenb[14]
port 293 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_oenb[15]
port 294 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oenb[16]
port 295 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[17]
port 296 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_oenb[18]
port 297 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_oenb[19]
port 298 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[1]
port 299 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_oenb[20]
port 300 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_oenb[21]
port 301 nsew signal input
rlabel metal2 s 165342 0 165398 800 6 la_oenb[22]
port 302 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_oenb[23]
port 303 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_oenb[24]
port 304 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 la_oenb[25]
port 305 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_oenb[26]
port 306 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oenb[27]
port 307 nsew signal input
rlabel metal2 s 180246 0 180302 800 6 la_oenb[28]
port 308 nsew signal input
rlabel metal2 s 182730 0 182786 800 6 la_oenb[29]
port 309 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_oenb[2]
port 310 nsew signal input
rlabel metal2 s 185214 0 185270 800 6 la_oenb[30]
port 311 nsew signal input
rlabel metal2 s 187698 0 187754 800 6 la_oenb[31]
port 312 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 la_oenb[32]
port 313 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 la_oenb[33]
port 314 nsew signal input
rlabel metal2 s 195150 0 195206 800 6 la_oenb[34]
port 315 nsew signal input
rlabel metal2 s 197634 0 197690 800 6 la_oenb[35]
port 316 nsew signal input
rlabel metal2 s 200118 0 200174 800 6 la_oenb[36]
port 317 nsew signal input
rlabel metal2 s 202602 0 202658 800 6 la_oenb[37]
port 318 nsew signal input
rlabel metal2 s 205086 0 205142 800 6 la_oenb[38]
port 319 nsew signal input
rlabel metal2 s 207570 0 207626 800 6 la_oenb[39]
port 320 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_oenb[3]
port 321 nsew signal input
rlabel metal2 s 210054 0 210110 800 6 la_oenb[40]
port 322 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_oenb[41]
port 323 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_oenb[42]
port 324 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_oenb[43]
port 325 nsew signal input
rlabel metal2 s 219990 0 220046 800 6 la_oenb[44]
port 326 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_oenb[45]
port 327 nsew signal input
rlabel metal2 s 224958 0 225014 800 6 la_oenb[46]
port 328 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 la_oenb[47]
port 329 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_oenb[48]
port 330 nsew signal input
rlabel metal2 s 232410 0 232466 800 6 la_oenb[49]
port 331 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_oenb[4]
port 332 nsew signal input
rlabel metal2 s 234894 0 234950 800 6 la_oenb[50]
port 333 nsew signal input
rlabel metal2 s 237378 0 237434 800 6 la_oenb[51]
port 334 nsew signal input
rlabel metal2 s 239862 0 239918 800 6 la_oenb[52]
port 335 nsew signal input
rlabel metal2 s 242346 0 242402 800 6 la_oenb[53]
port 336 nsew signal input
rlabel metal2 s 244830 0 244886 800 6 la_oenb[54]
port 337 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 la_oenb[55]
port 338 nsew signal input
rlabel metal2 s 249798 0 249854 800 6 la_oenb[56]
port 339 nsew signal input
rlabel metal2 s 252282 0 252338 800 6 la_oenb[57]
port 340 nsew signal input
rlabel metal2 s 254766 0 254822 800 6 la_oenb[58]
port 341 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_oenb[59]
port 342 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_oenb[5]
port 343 nsew signal input
rlabel metal2 s 259734 0 259790 800 6 la_oenb[60]
port 344 nsew signal input
rlabel metal2 s 262218 0 262274 800 6 la_oenb[61]
port 345 nsew signal input
rlabel metal2 s 264702 0 264758 800 6 la_oenb[62]
port 346 nsew signal input
rlabel metal2 s 267186 0 267242 800 6 la_oenb[63]
port 347 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 la_oenb[64]
port 348 nsew signal input
rlabel metal2 s 272154 0 272210 800 6 la_oenb[65]
port 349 nsew signal input
rlabel metal2 s 274638 0 274694 800 6 la_oenb[66]
port 350 nsew signal input
rlabel metal2 s 277122 0 277178 800 6 la_oenb[67]
port 351 nsew signal input
rlabel metal2 s 279606 0 279662 800 6 la_oenb[68]
port 352 nsew signal input
rlabel metal2 s 282090 0 282146 800 6 la_oenb[69]
port 353 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 la_oenb[6]
port 354 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 la_oenb[70]
port 355 nsew signal input
rlabel metal2 s 287058 0 287114 800 6 la_oenb[71]
port 356 nsew signal input
rlabel metal2 s 289542 0 289598 800 6 la_oenb[72]
port 357 nsew signal input
rlabel metal2 s 292026 0 292082 800 6 la_oenb[73]
port 358 nsew signal input
rlabel metal2 s 294510 0 294566 800 6 la_oenb[74]
port 359 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_oenb[75]
port 360 nsew signal input
rlabel metal2 s 299478 0 299534 800 6 la_oenb[76]
port 361 nsew signal input
rlabel metal2 s 301962 0 302018 800 6 la_oenb[77]
port 362 nsew signal input
rlabel metal2 s 304446 0 304502 800 6 la_oenb[78]
port 363 nsew signal input
rlabel metal2 s 306930 0 306986 800 6 la_oenb[79]
port 364 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oenb[7]
port 365 nsew signal input
rlabel metal2 s 309414 0 309470 800 6 la_oenb[80]
port 366 nsew signal input
rlabel metal2 s 311898 0 311954 800 6 la_oenb[81]
port 367 nsew signal input
rlabel metal2 s 314382 0 314438 800 6 la_oenb[82]
port 368 nsew signal input
rlabel metal2 s 316866 0 316922 800 6 la_oenb[83]
port 369 nsew signal input
rlabel metal2 s 319350 0 319406 800 6 la_oenb[84]
port 370 nsew signal input
rlabel metal2 s 321834 0 321890 800 6 la_oenb[85]
port 371 nsew signal input
rlabel metal2 s 324318 0 324374 800 6 la_oenb[86]
port 372 nsew signal input
rlabel metal2 s 326802 0 326858 800 6 la_oenb[87]
port 373 nsew signal input
rlabel metal2 s 329286 0 329342 800 6 la_oenb[88]
port 374 nsew signal input
rlabel metal2 s 331770 0 331826 800 6 la_oenb[89]
port 375 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_oenb[8]
port 376 nsew signal input
rlabel metal2 s 334254 0 334310 800 6 la_oenb[90]
port 377 nsew signal input
rlabel metal2 s 336738 0 336794 800 6 la_oenb[91]
port 378 nsew signal input
rlabel metal2 s 339222 0 339278 800 6 la_oenb[92]
port 379 nsew signal input
rlabel metal2 s 341706 0 341762 800 6 la_oenb[93]
port 380 nsew signal input
rlabel metal2 s 344190 0 344246 800 6 la_oenb[94]
port 381 nsew signal input
rlabel metal2 s 346674 0 346730 800 6 la_oenb[95]
port 382 nsew signal input
rlabel metal2 s 349158 0 349214 800 6 la_oenb[96]
port 383 nsew signal input
rlabel metal2 s 351642 0 351698 800 6 la_oenb[97]
port 384 nsew signal input
rlabel metal2 s 354126 0 354182 800 6 la_oenb[98]
port 385 nsew signal input
rlabel metal2 s 356610 0 356666 800 6 la_oenb[99]
port 386 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[9]
port 387 nsew signal input
rlabel metal4 s 4208 2128 4528 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 447760 6 vccd1
port 388 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 447760 6 vssd1
port 389 nsew ground bidirectional
rlabel metal2 s 21270 0 21326 800 6 wb_clk_i
port 390 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wb_rst_i
port 391 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_ack_o
port 392 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_adr_i[0]
port 393 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_adr_i[10]
port 394 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_adr_i[11]
port 395 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 wbs_adr_i[12]
port 396 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_adr_i[13]
port 397 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 wbs_adr_i[14]
port 398 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_adr_i[15]
port 399 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wbs_adr_i[16]
port 400 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 wbs_adr_i[17]
port 401 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 wbs_adr_i[18]
port 402 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 wbs_adr_i[19]
port 403 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[1]
port 404 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 wbs_adr_i[20]
port 405 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 wbs_adr_i[21]
port 406 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 wbs_adr_i[22]
port 407 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 wbs_adr_i[23]
port 408 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_adr_i[24]
port 409 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 wbs_adr_i[25]
port 410 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 wbs_adr_i[26]
port 411 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 wbs_adr_i[27]
port 412 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 wbs_adr_i[28]
port 413 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 wbs_adr_i[29]
port 414 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[2]
port 415 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 wbs_adr_i[30]
port 416 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 wbs_adr_i[31]
port 417 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_adr_i[3]
port 418 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[4]
port 419 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[5]
port 420 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_adr_i[6]
port 421 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_adr_i[7]
port 422 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_adr_i[8]
port 423 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_adr_i[9]
port 424 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_cyc_i
port 425 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_i[0]
port 426 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_i[10]
port 427 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_dat_i[11]
port 428 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 wbs_dat_i[12]
port 429 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 wbs_dat_i[13]
port 430 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 wbs_dat_i[14]
port 431 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_i[15]
port 432 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 wbs_dat_i[16]
port 433 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 wbs_dat_i[17]
port 434 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 wbs_dat_i[18]
port 435 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_i[19]
port 436 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_i[1]
port 437 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 wbs_dat_i[20]
port 438 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 wbs_dat_i[21]
port 439 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 wbs_dat_i[22]
port 440 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 wbs_dat_i[23]
port 441 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 wbs_dat_i[24]
port 442 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_i[25]
port 443 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 wbs_dat_i[26]
port 444 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 wbs_dat_i[27]
port 445 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 wbs_dat_i[28]
port 446 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 wbs_dat_i[29]
port 447 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[2]
port 448 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 wbs_dat_i[30]
port 449 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 wbs_dat_i[31]
port 450 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_i[3]
port 451 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_i[4]
port 452 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[5]
port 453 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_i[6]
port 454 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 wbs_dat_i[7]
port 455 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_i[8]
port 456 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_dat_i[9]
port 457 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[0]
port 458 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 wbs_dat_o[10]
port 459 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 wbs_dat_o[11]
port 460 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 wbs_dat_o[12]
port 461 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 wbs_dat_o[13]
port 462 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 wbs_dat_o[14]
port 463 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 wbs_dat_o[15]
port 464 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_o[16]
port 465 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 wbs_dat_o[17]
port 466 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 wbs_dat_o[18]
port 467 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 wbs_dat_o[19]
port 468 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[1]
port 469 nsew signal output
rlabel metal2 s 80886 0 80942 800 6 wbs_dat_o[20]
port 470 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 wbs_dat_o[21]
port 471 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 wbs_dat_o[22]
port 472 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 wbs_dat_o[23]
port 473 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 wbs_dat_o[24]
port 474 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 wbs_dat_o[25]
port 475 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 wbs_dat_o[26]
port 476 nsew signal output
rlabel metal2 s 98274 0 98330 800 6 wbs_dat_o[27]
port 477 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 wbs_dat_o[28]
port 478 nsew signal output
rlabel metal2 s 103242 0 103298 800 6 wbs_dat_o[29]
port 479 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_o[2]
port 480 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 wbs_dat_o[30]
port 481 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 wbs_dat_o[31]
port 482 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_o[3]
port 483 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[4]
port 484 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_o[5]
port 485 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_o[6]
port 486 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[7]
port 487 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_o[8]
port 488 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 wbs_dat_o[9]
port 489 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_sel_i[0]
port 490 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 wbs_sel_i[1]
port 491 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_sel_i[2]
port 492 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_sel_i[3]
port 493 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_stb_i
port 494 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_we_i
port 495 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 450000 450000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 65321924
string GDS_FILE /home/wouter/openmpw/caravel_labs_search/openlane/user_proj_example/runs/22_08_13_14_46/results/signoff/user_proj_example.magic.gds
string GDS_START 1001478
<< end >>

