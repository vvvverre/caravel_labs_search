VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2250.000 BY 2250.000 ;
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2134.950 0.000 2135.230 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2139.090 0.000 2139.370 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.230 0.000 2143.510 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 0.000 1787.470 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.610 0.000 1799.890 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.030 0.000 1812.310 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.450 0.000 1824.730 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1836.870 0.000 1837.150 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.290 0.000 1849.570 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.710 0.000 1861.990 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.130 0.000 1874.410 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.550 0.000 1886.830 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.970 0.000 1899.250 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 0.000 669.670 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.390 0.000 1911.670 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.810 0.000 1924.090 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.230 0.000 1936.510 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.650 0.000 1948.930 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.070 0.000 1961.350 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.490 0.000 1973.770 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.910 0.000 1986.190 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.330 0.000 1998.610 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2010.750 0.000 2011.030 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.170 0.000 2023.450 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.590 0.000 2035.870 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.010 0.000 2048.290 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.430 0.000 2060.710 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2072.850 0.000 2073.130 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.270 0.000 2085.550 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2097.690 0.000 2097.970 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2110.110 0.000 2110.390 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.530 0.000 2122.810 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 0.000 706.930 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.330 0.000 756.610 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 0.000 868.390 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.530 0.000 880.810 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 0.000 893.230 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 0.000 905.650 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 0.000 930.490 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.630 0.000 942.910 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 0.000 955.330 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 0.000 980.170 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 0.000 992.590 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.150 0.000 1017.430 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.990 0.000 1042.270 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 0.000 1054.690 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.830 0.000 1067.110 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 0.000 1079.530 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 0.000 1091.950 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 0.000 1116.790 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.930 0.000 1129.210 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.350 0.000 1141.630 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.770 0.000 1154.050 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.190 0.000 1166.470 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.030 0.000 1191.310 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.450 0.000 1203.730 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1215.870 0.000 1216.150 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.290 0.000 1228.570 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.710 0.000 1240.990 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 0.000 1253.410 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1277.970 0.000 1278.250 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.390 0.000 1290.670 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.810 0.000 1303.090 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.230 0.000 1315.510 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.650 0.000 1327.930 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.070 0.000 1340.350 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1364.910 0.000 1365.190 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1377.330 0.000 1377.610 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.750 0.000 1390.030 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1402.170 0.000 1402.450 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.590 0.000 1414.870 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1427.010 0.000 1427.290 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 0.000 1439.710 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.850 0.000 1452.130 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.270 0.000 1464.550 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1476.690 0.000 1476.970 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 0.000 1489.390 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1501.530 0.000 1501.810 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.950 0.000 1514.230 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 0.000 1526.650 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1538.790 0.000 1539.070 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.210 0.000 1551.490 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.630 0.000 1563.910 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.050 0.000 1576.330 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.470 0.000 1588.750 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.890 0.000 1601.170 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.310 0.000 1613.590 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 0.000 1626.010 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.150 0.000 1638.430 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.570 0.000 1650.850 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.990 0.000 1663.270 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.410 0.000 1675.690 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.830 0.000 1688.110 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1700.250 0.000 1700.530 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.670 0.000 1712.950 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.090 0.000 1725.370 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.510 0.000 1737.790 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.930 0.000 1750.210 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.350 0.000 1762.630 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1774.770 0.000 1775.050 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1791.330 0.000 1791.610 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.750 0.000 1804.030 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 0.000 1816.450 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.590 0.000 1828.870 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.010 0.000 1841.290 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.430 0.000 1853.710 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.850 0.000 1866.130 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.270 0.000 1878.550 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.690 0.000 1890.970 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.110 0.000 1903.390 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 0.000 673.810 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.530 0.000 1915.810 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.950 0.000 1928.230 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.370 0.000 1940.650 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1952.790 0.000 1953.070 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.210 0.000 1965.490 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.630 0.000 1977.910 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.050 0.000 1990.330 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.470 0.000 2002.750 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.890 0.000 2015.170 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.310 0.000 2027.590 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.730 0.000 2040.010 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.150 0.000 2052.430 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.570 0.000 2064.850 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2076.990 0.000 2077.270 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.410 0.000 2089.690 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2101.830 0.000 2102.110 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2114.250 0.000 2114.530 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.670 0.000 2126.950 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 0.000 835.270 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.410 0.000 847.690 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 0.000 860.110 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 0.000 872.530 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.670 0.000 884.950 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 0.000 897.370 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.930 0.000 922.210 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 0.000 934.630 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.770 0.000 947.050 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 0.000 959.470 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.610 0.000 971.890 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.030 0.000 984.310 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 0.000 996.730 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1008.870 0.000 1009.150 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 0.000 1021.570 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.710 0.000 1033.990 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 0.000 1058.830 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.970 0.000 1071.250 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.390 0.000 1083.670 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 0.000 1096.090 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.230 0.000 1108.510 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.650 0.000 1120.930 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.070 0.000 1133.350 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 0.000 1145.770 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.910 0.000 1158.190 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.330 0.000 1170.610 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.750 0.000 1183.030 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.010 0.000 1220.290 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.430 0.000 1232.710 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1244.850 0.000 1245.130 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 0.000 1257.550 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 0.000 1269.970 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.110 0.000 1282.390 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.530 0.000 1294.810 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1306.950 0.000 1307.230 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 0.000 1319.650 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.790 0.000 1332.070 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 0.000 1344.490 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.630 0.000 1356.910 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.050 0.000 1369.330 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.470 0.000 1381.750 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.890 0.000 1394.170 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.310 0.000 1406.590 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 0.000 1419.010 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.150 0.000 1431.430 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1443.570 0.000 1443.850 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 0.000 1456.270 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.830 0.000 1481.110 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1493.250 0.000 1493.530 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1505.670 0.000 1505.950 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.090 0.000 1518.370 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.510 0.000 1530.790 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 0.000 1543.210 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 0.000 1555.630 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.770 0.000 1568.050 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.190 0.000 1580.470 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.610 0.000 1592.890 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.030 0.000 1605.310 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.450 0.000 1617.730 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1629.870 0.000 1630.150 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1642.290 0.000 1642.570 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.710 0.000 1654.990 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.130 0.000 1667.410 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.550 0.000 1679.830 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 0.000 1692.250 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.390 0.000 1704.670 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.810 0.000 1717.090 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.230 0.000 1729.510 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.650 0.000 1741.930 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.070 0.000 1754.350 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.490 0.000 1766.770 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1778.910 0.000 1779.190 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 0.000 553.750 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.470 0.000 1795.750 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1807.890 0.000 1808.170 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1820.310 0.000 1820.590 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.730 0.000 1833.010 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.150 0.000 1845.430 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.570 0.000 1857.850 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.990 0.000 1870.270 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.410 0.000 1882.690 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.830 0.000 1895.110 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1907.250 0.000 1907.530 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.670 0.000 1919.950 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.090 0.000 1932.370 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.510 0.000 1944.790 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.930 0.000 1957.210 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.350 0.000 1969.630 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.770 0.000 1982.050 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.190 0.000 1994.470 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.610 0.000 2006.890 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.030 0.000 2019.310 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2031.450 0.000 2031.730 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2043.870 0.000 2044.150 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2056.290 0.000 2056.570 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.710 0.000 2068.990 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2081.130 0.000 2081.410 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.550 0.000 2093.830 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.970 0.000 2106.250 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.390 0.000 2118.670 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.810 0.000 2131.090 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 0.000 826.990 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 0.000 839.410 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.550 0.000 851.830 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.970 0.000 864.250 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 0.000 926.350 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 0.000 938.770 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 0.000 963.610 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.750 0.000 976.030 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.170 0.000 988.450 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.430 0.000 1025.710 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.850 0.000 1038.130 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 0.000 1050.550 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.110 0.000 1075.390 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 0.000 1087.810 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 0.000 1100.230 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1112.370 0.000 1112.650 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 0.000 1125.070 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 0.000 1162.330 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 0.000 603.430 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.470 0.000 1174.750 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 0.000 1187.170 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.310 0.000 1199.590 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.730 0.000 1212.010 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 0.000 1224.430 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1236.570 0.000 1236.850 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1248.990 0.000 1249.270 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.410 0.000 1261.690 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 0.000 1274.110 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.250 0.000 1286.530 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.670 0.000 1298.950 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.090 0.000 1311.370 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 0.000 1323.790 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.930 0.000 1336.210 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 0.000 1361.050 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.190 0.000 1373.470 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.610 0.000 1385.890 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.030 0.000 1398.310 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 0.000 1435.570 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1447.710 0.000 1447.990 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.130 0.000 1460.410 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.550 0.000 1472.830 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.970 0.000 1485.250 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 0.000 1497.670 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.810 0.000 1510.090 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.230 0.000 1522.510 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.650 0.000 1534.930 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.070 0.000 1547.350 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.490 0.000 1559.770 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.910 0.000 1572.190 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.330 0.000 1584.610 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.750 0.000 1597.030 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.170 0.000 1609.450 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.590 0.000 1621.870 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.010 0.000 1634.290 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.430 0.000 1646.710 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.850 0.000 1659.130 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 0.000 653.110 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.270 0.000 1671.550 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.690 0.000 1683.970 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.110 0.000 1696.390 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.530 0.000 1708.810 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.950 0.000 1721.230 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1733.370 0.000 1733.650 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.790 0.000 1746.070 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.210 0.000 1758.490 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.630 0.000 1770.910 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.050 0.000 1783.330 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 2238.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 2238.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 2238.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 0.000 321.910 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 0.000 247.390 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 0.000 450.250 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 0.000 239.110 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 0.000 429.550 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.210 0.000 516.490 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER nwell ;
        RECT 5.330 2237.145 2244.530 2238.750 ;
        RECT 5.330 2231.705 2244.530 2234.535 ;
        RECT 5.330 2226.265 2244.530 2229.095 ;
        RECT 5.330 2220.825 2244.530 2223.655 ;
        RECT 5.330 2215.385 2244.530 2218.215 ;
        RECT 5.330 2209.945 2244.530 2212.775 ;
        RECT 5.330 2204.505 2244.530 2207.335 ;
        RECT 5.330 2199.065 2244.530 2201.895 ;
        RECT 5.330 2193.625 2244.530 2196.455 ;
        RECT 5.330 2188.185 2244.530 2191.015 ;
        RECT 5.330 2182.745 2244.530 2185.575 ;
        RECT 5.330 2177.305 2244.530 2180.135 ;
        RECT 5.330 2171.865 2244.530 2174.695 ;
        RECT 5.330 2166.425 2244.530 2169.255 ;
        RECT 5.330 2160.985 2244.530 2163.815 ;
        RECT 5.330 2155.545 2244.530 2158.375 ;
        RECT 5.330 2150.105 2244.530 2152.935 ;
        RECT 5.330 2144.665 2244.530 2147.495 ;
        RECT 5.330 2139.225 2244.530 2142.055 ;
        RECT 5.330 2133.785 2244.530 2136.615 ;
        RECT 5.330 2128.345 2244.530 2131.175 ;
        RECT 5.330 2122.905 2244.530 2125.735 ;
        RECT 5.330 2117.465 2244.530 2120.295 ;
        RECT 5.330 2112.025 2244.530 2114.855 ;
        RECT 5.330 2106.585 2244.530 2109.415 ;
        RECT 5.330 2101.145 2244.530 2103.975 ;
        RECT 5.330 2095.705 2244.530 2098.535 ;
        RECT 5.330 2090.265 2244.530 2093.095 ;
        RECT 5.330 2084.825 2244.530 2087.655 ;
        RECT 5.330 2079.385 2244.530 2082.215 ;
        RECT 5.330 2073.945 2244.530 2076.775 ;
        RECT 5.330 2068.505 2244.530 2071.335 ;
        RECT 5.330 2063.065 2244.530 2065.895 ;
        RECT 5.330 2057.625 2244.530 2060.455 ;
        RECT 5.330 2052.185 2244.530 2055.015 ;
        RECT 5.330 2046.745 2244.530 2049.575 ;
        RECT 5.330 2041.305 2244.530 2044.135 ;
        RECT 5.330 2035.865 2244.530 2038.695 ;
        RECT 5.330 2030.425 2244.530 2033.255 ;
        RECT 5.330 2024.985 2244.530 2027.815 ;
        RECT 5.330 2019.545 2244.530 2022.375 ;
        RECT 5.330 2014.105 2244.530 2016.935 ;
        RECT 5.330 2008.665 2244.530 2011.495 ;
        RECT 5.330 2003.225 2244.530 2006.055 ;
        RECT 5.330 1997.785 2244.530 2000.615 ;
        RECT 5.330 1992.345 2244.530 1995.175 ;
        RECT 5.330 1986.905 2244.530 1989.735 ;
        RECT 5.330 1981.465 2244.530 1984.295 ;
        RECT 5.330 1976.025 2244.530 1978.855 ;
        RECT 5.330 1970.585 2244.530 1973.415 ;
        RECT 5.330 1965.145 2244.530 1967.975 ;
        RECT 5.330 1959.705 2244.530 1962.535 ;
        RECT 5.330 1954.265 2244.530 1957.095 ;
        RECT 5.330 1948.825 2244.530 1951.655 ;
        RECT 5.330 1943.385 2244.530 1946.215 ;
        RECT 5.330 1937.945 2244.530 1940.775 ;
        RECT 5.330 1932.505 2244.530 1935.335 ;
        RECT 5.330 1927.065 2244.530 1929.895 ;
        RECT 5.330 1921.625 2244.530 1924.455 ;
        RECT 5.330 1916.185 2244.530 1919.015 ;
        RECT 5.330 1910.745 2244.530 1913.575 ;
        RECT 5.330 1905.305 2244.530 1908.135 ;
        RECT 5.330 1899.865 2244.530 1902.695 ;
        RECT 5.330 1894.425 2244.530 1897.255 ;
        RECT 5.330 1888.985 2244.530 1891.815 ;
        RECT 5.330 1883.545 2244.530 1886.375 ;
        RECT 5.330 1878.105 2244.530 1880.935 ;
        RECT 5.330 1872.665 2244.530 1875.495 ;
        RECT 5.330 1867.225 2244.530 1870.055 ;
        RECT 5.330 1861.785 2244.530 1864.615 ;
        RECT 5.330 1856.345 2244.530 1859.175 ;
        RECT 5.330 1850.905 2244.530 1853.735 ;
        RECT 5.330 1845.465 2244.530 1848.295 ;
        RECT 5.330 1840.025 2244.530 1842.855 ;
        RECT 5.330 1834.585 2244.530 1837.415 ;
        RECT 5.330 1829.145 2244.530 1831.975 ;
        RECT 5.330 1823.705 2244.530 1826.535 ;
        RECT 5.330 1818.265 2244.530 1821.095 ;
        RECT 5.330 1812.825 2244.530 1815.655 ;
        RECT 5.330 1807.385 2244.530 1810.215 ;
        RECT 5.330 1801.945 2244.530 1804.775 ;
        RECT 5.330 1796.505 2244.530 1799.335 ;
        RECT 5.330 1791.065 2244.530 1793.895 ;
        RECT 5.330 1785.625 2244.530 1788.455 ;
        RECT 5.330 1780.185 2244.530 1783.015 ;
        RECT 5.330 1774.745 2244.530 1777.575 ;
        RECT 5.330 1769.305 2244.530 1772.135 ;
        RECT 5.330 1763.865 2244.530 1766.695 ;
        RECT 5.330 1758.425 2244.530 1761.255 ;
        RECT 5.330 1752.985 2244.530 1755.815 ;
        RECT 5.330 1747.545 2244.530 1750.375 ;
        RECT 5.330 1742.105 2244.530 1744.935 ;
        RECT 5.330 1736.665 2244.530 1739.495 ;
        RECT 5.330 1731.225 2244.530 1734.055 ;
        RECT 5.330 1725.785 2244.530 1728.615 ;
        RECT 5.330 1720.345 2244.530 1723.175 ;
        RECT 5.330 1714.905 2244.530 1717.735 ;
        RECT 5.330 1709.465 2244.530 1712.295 ;
        RECT 5.330 1704.025 2244.530 1706.855 ;
        RECT 5.330 1698.585 2244.530 1701.415 ;
        RECT 5.330 1693.145 2244.530 1695.975 ;
        RECT 5.330 1687.705 2244.530 1690.535 ;
        RECT 5.330 1682.265 2244.530 1685.095 ;
        RECT 5.330 1676.825 2244.530 1679.655 ;
        RECT 5.330 1671.385 2244.530 1674.215 ;
        RECT 5.330 1665.945 2244.530 1668.775 ;
        RECT 5.330 1660.505 2244.530 1663.335 ;
        RECT 5.330 1655.065 2244.530 1657.895 ;
        RECT 5.330 1649.625 2244.530 1652.455 ;
        RECT 5.330 1644.185 2244.530 1647.015 ;
        RECT 5.330 1638.745 2244.530 1641.575 ;
        RECT 5.330 1633.305 2244.530 1636.135 ;
        RECT 5.330 1627.865 2244.530 1630.695 ;
        RECT 5.330 1622.425 2244.530 1625.255 ;
        RECT 5.330 1616.985 2244.530 1619.815 ;
        RECT 5.330 1611.545 2244.530 1614.375 ;
        RECT 5.330 1606.105 2244.530 1608.935 ;
        RECT 5.330 1600.665 2244.530 1603.495 ;
        RECT 5.330 1595.225 2244.530 1598.055 ;
        RECT 5.330 1589.785 2244.530 1592.615 ;
        RECT 5.330 1584.345 2244.530 1587.175 ;
        RECT 5.330 1578.905 2244.530 1581.735 ;
        RECT 5.330 1573.465 2244.530 1576.295 ;
        RECT 5.330 1568.025 2244.530 1570.855 ;
        RECT 5.330 1562.585 2244.530 1565.415 ;
        RECT 5.330 1557.145 2244.530 1559.975 ;
        RECT 5.330 1551.705 2244.530 1554.535 ;
        RECT 5.330 1546.265 2244.530 1549.095 ;
        RECT 5.330 1540.825 2244.530 1543.655 ;
        RECT 5.330 1535.385 2244.530 1538.215 ;
        RECT 5.330 1529.945 2244.530 1532.775 ;
        RECT 5.330 1524.505 2244.530 1527.335 ;
        RECT 5.330 1519.065 2244.530 1521.895 ;
        RECT 5.330 1513.625 2244.530 1516.455 ;
        RECT 5.330 1508.185 2244.530 1511.015 ;
        RECT 5.330 1502.745 2244.530 1505.575 ;
        RECT 5.330 1497.305 2244.530 1500.135 ;
        RECT 5.330 1491.865 2244.530 1494.695 ;
        RECT 5.330 1486.425 2244.530 1489.255 ;
        RECT 5.330 1480.985 2244.530 1483.815 ;
        RECT 5.330 1475.545 2244.530 1478.375 ;
        RECT 5.330 1470.105 2244.530 1472.935 ;
        RECT 5.330 1464.665 2244.530 1467.495 ;
        RECT 5.330 1459.225 2244.530 1462.055 ;
        RECT 5.330 1453.785 2244.530 1456.615 ;
        RECT 5.330 1448.345 2244.530 1451.175 ;
        RECT 5.330 1442.905 2244.530 1445.735 ;
        RECT 5.330 1437.465 2244.530 1440.295 ;
        RECT 5.330 1432.025 2244.530 1434.855 ;
        RECT 5.330 1426.585 2244.530 1429.415 ;
        RECT 5.330 1421.145 2244.530 1423.975 ;
        RECT 5.330 1415.705 2244.530 1418.535 ;
        RECT 5.330 1410.265 2244.530 1413.095 ;
        RECT 5.330 1404.825 2244.530 1407.655 ;
        RECT 5.330 1399.385 2244.530 1402.215 ;
        RECT 5.330 1393.945 2244.530 1396.775 ;
        RECT 5.330 1388.505 2244.530 1391.335 ;
        RECT 5.330 1383.065 2244.530 1385.895 ;
        RECT 5.330 1377.625 2244.530 1380.455 ;
        RECT 5.330 1372.185 2244.530 1375.015 ;
        RECT 5.330 1366.745 2244.530 1369.575 ;
        RECT 5.330 1361.305 2244.530 1364.135 ;
        RECT 5.330 1355.865 2244.530 1358.695 ;
        RECT 5.330 1350.425 2244.530 1353.255 ;
        RECT 5.330 1344.985 2244.530 1347.815 ;
        RECT 5.330 1339.545 2244.530 1342.375 ;
        RECT 5.330 1334.105 2244.530 1336.935 ;
        RECT 5.330 1328.665 2244.530 1331.495 ;
        RECT 5.330 1323.225 2244.530 1326.055 ;
        RECT 5.330 1317.785 2244.530 1320.615 ;
        RECT 5.330 1312.345 2244.530 1315.175 ;
        RECT 5.330 1306.905 2244.530 1309.735 ;
        RECT 5.330 1301.465 2244.530 1304.295 ;
        RECT 5.330 1296.025 2244.530 1298.855 ;
        RECT 5.330 1290.585 2244.530 1293.415 ;
        RECT 5.330 1285.145 2244.530 1287.975 ;
        RECT 5.330 1279.705 2244.530 1282.535 ;
        RECT 5.330 1274.265 2244.530 1277.095 ;
        RECT 5.330 1268.825 2244.530 1271.655 ;
        RECT 5.330 1263.385 2244.530 1266.215 ;
        RECT 5.330 1257.945 2244.530 1260.775 ;
        RECT 5.330 1252.505 2244.530 1255.335 ;
        RECT 5.330 1247.065 2244.530 1249.895 ;
        RECT 5.330 1241.625 2244.530 1244.455 ;
        RECT 5.330 1236.185 2244.530 1239.015 ;
        RECT 5.330 1230.745 2244.530 1233.575 ;
        RECT 5.330 1225.305 2244.530 1228.135 ;
        RECT 5.330 1219.865 2244.530 1222.695 ;
        RECT 5.330 1214.425 2244.530 1217.255 ;
        RECT 5.330 1208.985 2244.530 1211.815 ;
        RECT 5.330 1203.545 2244.530 1206.375 ;
        RECT 5.330 1198.105 2244.530 1200.935 ;
        RECT 5.330 1192.665 2244.530 1195.495 ;
        RECT 5.330 1187.225 2244.530 1190.055 ;
        RECT 5.330 1181.785 2244.530 1184.615 ;
        RECT 5.330 1176.345 2244.530 1179.175 ;
        RECT 5.330 1170.905 2244.530 1173.735 ;
        RECT 5.330 1165.465 2244.530 1168.295 ;
        RECT 5.330 1160.025 2244.530 1162.855 ;
        RECT 5.330 1154.585 2244.530 1157.415 ;
        RECT 5.330 1149.145 2244.530 1151.975 ;
        RECT 5.330 1143.705 2244.530 1146.535 ;
        RECT 5.330 1138.265 2244.530 1141.095 ;
        RECT 5.330 1132.825 2244.530 1135.655 ;
        RECT 5.330 1127.385 2244.530 1130.215 ;
        RECT 5.330 1121.945 2244.530 1124.775 ;
        RECT 5.330 1116.505 2244.530 1119.335 ;
        RECT 5.330 1111.065 2244.530 1113.895 ;
        RECT 5.330 1105.625 2244.530 1108.455 ;
        RECT 5.330 1100.185 2244.530 1103.015 ;
        RECT 5.330 1094.745 2244.530 1097.575 ;
        RECT 5.330 1089.305 2244.530 1092.135 ;
        RECT 5.330 1083.865 2244.530 1086.695 ;
        RECT 5.330 1078.425 2244.530 1081.255 ;
        RECT 5.330 1072.985 2244.530 1075.815 ;
        RECT 5.330 1067.545 2244.530 1070.375 ;
        RECT 5.330 1062.105 2244.530 1064.935 ;
        RECT 5.330 1056.665 2244.530 1059.495 ;
        RECT 5.330 1051.225 2244.530 1054.055 ;
        RECT 5.330 1045.785 2244.530 1048.615 ;
        RECT 5.330 1040.345 2244.530 1043.175 ;
        RECT 5.330 1034.905 2244.530 1037.735 ;
        RECT 5.330 1029.465 2244.530 1032.295 ;
        RECT 5.330 1024.025 2244.530 1026.855 ;
        RECT 5.330 1018.585 2244.530 1021.415 ;
        RECT 5.330 1013.145 2244.530 1015.975 ;
        RECT 5.330 1007.705 2244.530 1010.535 ;
        RECT 5.330 1002.265 2244.530 1005.095 ;
        RECT 5.330 996.825 2244.530 999.655 ;
        RECT 5.330 991.385 2244.530 994.215 ;
        RECT 5.330 985.945 2244.530 988.775 ;
        RECT 5.330 980.505 2244.530 983.335 ;
        RECT 5.330 975.065 2244.530 977.895 ;
        RECT 5.330 969.625 2244.530 972.455 ;
        RECT 5.330 964.185 2244.530 967.015 ;
        RECT 5.330 958.745 2244.530 961.575 ;
        RECT 5.330 953.305 2244.530 956.135 ;
        RECT 5.330 947.865 2244.530 950.695 ;
        RECT 5.330 942.425 2244.530 945.255 ;
        RECT 5.330 936.985 2244.530 939.815 ;
        RECT 5.330 931.545 2244.530 934.375 ;
        RECT 5.330 926.105 2244.530 928.935 ;
        RECT 5.330 920.665 2244.530 923.495 ;
        RECT 5.330 915.225 2244.530 918.055 ;
        RECT 5.330 909.785 2244.530 912.615 ;
        RECT 5.330 904.345 2244.530 907.175 ;
        RECT 5.330 898.905 2244.530 901.735 ;
        RECT 5.330 893.465 2244.530 896.295 ;
        RECT 5.330 888.025 2244.530 890.855 ;
        RECT 5.330 882.585 2244.530 885.415 ;
        RECT 5.330 877.145 2244.530 879.975 ;
        RECT 5.330 871.705 2244.530 874.535 ;
        RECT 5.330 866.265 2244.530 869.095 ;
        RECT 5.330 860.825 2244.530 863.655 ;
        RECT 5.330 855.385 2244.530 858.215 ;
        RECT 5.330 849.945 2244.530 852.775 ;
        RECT 5.330 844.505 2244.530 847.335 ;
        RECT 5.330 839.065 2244.530 841.895 ;
        RECT 5.330 833.625 2244.530 836.455 ;
        RECT 5.330 828.185 2244.530 831.015 ;
        RECT 5.330 822.745 2244.530 825.575 ;
        RECT 5.330 817.305 2244.530 820.135 ;
        RECT 5.330 811.865 2244.530 814.695 ;
        RECT 5.330 806.425 2244.530 809.255 ;
        RECT 5.330 800.985 2244.530 803.815 ;
        RECT 5.330 795.545 2244.530 798.375 ;
        RECT 5.330 790.105 2244.530 792.935 ;
        RECT 5.330 784.665 2244.530 787.495 ;
        RECT 5.330 779.225 2244.530 782.055 ;
        RECT 5.330 773.785 2244.530 776.615 ;
        RECT 5.330 768.345 2244.530 771.175 ;
        RECT 5.330 762.905 2244.530 765.735 ;
        RECT 5.330 757.465 2244.530 760.295 ;
        RECT 5.330 752.025 2244.530 754.855 ;
        RECT 5.330 746.585 2244.530 749.415 ;
        RECT 5.330 741.145 2244.530 743.975 ;
        RECT 5.330 735.705 2244.530 738.535 ;
        RECT 5.330 730.265 2244.530 733.095 ;
        RECT 5.330 724.825 2244.530 727.655 ;
        RECT 5.330 719.385 2244.530 722.215 ;
        RECT 5.330 713.945 2244.530 716.775 ;
        RECT 5.330 708.505 2244.530 711.335 ;
        RECT 5.330 703.065 2244.530 705.895 ;
        RECT 5.330 697.625 2244.530 700.455 ;
        RECT 5.330 692.185 2244.530 695.015 ;
        RECT 5.330 686.745 2244.530 689.575 ;
        RECT 5.330 681.305 2244.530 684.135 ;
        RECT 5.330 675.865 2244.530 678.695 ;
        RECT 5.330 670.425 2244.530 673.255 ;
        RECT 5.330 664.985 2244.530 667.815 ;
        RECT 5.330 659.545 2244.530 662.375 ;
        RECT 5.330 654.105 2244.530 656.935 ;
        RECT 5.330 648.665 2244.530 651.495 ;
        RECT 5.330 643.225 2244.530 646.055 ;
        RECT 5.330 637.785 2244.530 640.615 ;
        RECT 5.330 632.345 2244.530 635.175 ;
        RECT 5.330 626.905 2244.530 629.735 ;
        RECT 5.330 621.465 2244.530 624.295 ;
        RECT 5.330 616.025 2244.530 618.855 ;
        RECT 5.330 610.585 2244.530 613.415 ;
        RECT 5.330 605.145 2244.530 607.975 ;
        RECT 5.330 599.705 2244.530 602.535 ;
        RECT 5.330 594.265 2244.530 597.095 ;
        RECT 5.330 588.825 2244.530 591.655 ;
        RECT 5.330 583.385 2244.530 586.215 ;
        RECT 5.330 577.945 2244.530 580.775 ;
        RECT 5.330 572.505 2244.530 575.335 ;
        RECT 5.330 567.065 2244.530 569.895 ;
        RECT 5.330 561.625 2244.530 564.455 ;
        RECT 5.330 556.185 2244.530 559.015 ;
        RECT 5.330 550.745 2244.530 553.575 ;
        RECT 5.330 545.305 2244.530 548.135 ;
        RECT 5.330 539.865 2244.530 542.695 ;
        RECT 5.330 534.425 2244.530 537.255 ;
        RECT 5.330 528.985 2244.530 531.815 ;
        RECT 5.330 523.545 2244.530 526.375 ;
        RECT 5.330 518.105 2244.530 520.935 ;
        RECT 5.330 512.665 2244.530 515.495 ;
        RECT 5.330 507.225 2244.530 510.055 ;
        RECT 5.330 501.785 2244.530 504.615 ;
        RECT 5.330 496.345 2244.530 499.175 ;
        RECT 5.330 490.905 2244.530 493.735 ;
        RECT 5.330 485.465 2244.530 488.295 ;
        RECT 5.330 480.025 2244.530 482.855 ;
        RECT 5.330 474.585 2244.530 477.415 ;
        RECT 5.330 469.145 2244.530 471.975 ;
        RECT 5.330 463.705 2244.530 466.535 ;
        RECT 5.330 458.265 2244.530 461.095 ;
        RECT 5.330 452.825 2244.530 455.655 ;
        RECT 5.330 447.385 2244.530 450.215 ;
        RECT 5.330 441.945 2244.530 444.775 ;
        RECT 5.330 436.505 2244.530 439.335 ;
        RECT 5.330 431.065 2244.530 433.895 ;
        RECT 5.330 425.625 2244.530 428.455 ;
        RECT 5.330 420.185 2244.530 423.015 ;
        RECT 5.330 414.745 2244.530 417.575 ;
        RECT 5.330 409.305 2244.530 412.135 ;
        RECT 5.330 403.865 2244.530 406.695 ;
        RECT 5.330 398.425 2244.530 401.255 ;
        RECT 5.330 392.985 2244.530 395.815 ;
        RECT 5.330 387.545 2244.530 390.375 ;
        RECT 5.330 382.105 2244.530 384.935 ;
        RECT 5.330 376.665 2244.530 379.495 ;
        RECT 5.330 371.225 2244.530 374.055 ;
        RECT 5.330 365.785 2244.530 368.615 ;
        RECT 5.330 360.345 2244.530 363.175 ;
        RECT 5.330 354.905 2244.530 357.735 ;
        RECT 5.330 349.465 2244.530 352.295 ;
        RECT 5.330 344.025 2244.530 346.855 ;
        RECT 5.330 338.585 2244.530 341.415 ;
        RECT 5.330 333.145 2244.530 335.975 ;
        RECT 5.330 327.705 2244.530 330.535 ;
        RECT 5.330 322.265 2244.530 325.095 ;
        RECT 5.330 316.825 2244.530 319.655 ;
        RECT 5.330 311.385 2244.530 314.215 ;
        RECT 5.330 305.945 2244.530 308.775 ;
        RECT 5.330 300.505 2244.530 303.335 ;
        RECT 5.330 295.065 2244.530 297.895 ;
        RECT 5.330 289.625 2244.530 292.455 ;
        RECT 5.330 284.185 2244.530 287.015 ;
        RECT 5.330 278.745 2244.530 281.575 ;
        RECT 5.330 273.305 2244.530 276.135 ;
        RECT 5.330 267.865 2244.530 270.695 ;
        RECT 5.330 262.425 2244.530 265.255 ;
        RECT 5.330 256.985 2244.530 259.815 ;
        RECT 5.330 251.545 2244.530 254.375 ;
        RECT 5.330 246.105 2244.530 248.935 ;
        RECT 5.330 240.665 2244.530 243.495 ;
        RECT 5.330 235.225 2244.530 238.055 ;
        RECT 5.330 229.785 2244.530 232.615 ;
        RECT 5.330 224.345 2244.530 227.175 ;
        RECT 5.330 218.905 2244.530 221.735 ;
        RECT 5.330 213.465 2244.530 216.295 ;
        RECT 5.330 208.025 2244.530 210.855 ;
        RECT 5.330 202.585 2244.530 205.415 ;
        RECT 5.330 197.145 2244.530 199.975 ;
        RECT 5.330 191.705 2244.530 194.535 ;
        RECT 5.330 186.265 2244.530 189.095 ;
        RECT 5.330 180.825 2244.530 183.655 ;
        RECT 5.330 175.385 2244.530 178.215 ;
        RECT 5.330 169.945 2244.530 172.775 ;
        RECT 5.330 164.505 2244.530 167.335 ;
        RECT 5.330 159.065 2244.530 161.895 ;
        RECT 5.330 153.625 2244.530 156.455 ;
        RECT 5.330 148.185 2244.530 151.015 ;
        RECT 5.330 142.745 2244.530 145.575 ;
        RECT 5.330 137.305 2244.530 140.135 ;
        RECT 5.330 131.865 2244.530 134.695 ;
        RECT 5.330 126.425 2244.530 129.255 ;
        RECT 5.330 120.985 2244.530 123.815 ;
        RECT 5.330 115.545 2244.530 118.375 ;
        RECT 5.330 110.105 2244.530 112.935 ;
        RECT 5.330 104.665 2244.530 107.495 ;
        RECT 5.330 99.225 2244.530 102.055 ;
        RECT 5.330 93.785 2244.530 96.615 ;
        RECT 5.330 88.345 2244.530 91.175 ;
        RECT 5.330 82.905 2244.530 85.735 ;
        RECT 5.330 77.465 2244.530 80.295 ;
        RECT 5.330 72.025 2244.530 74.855 ;
        RECT 5.330 66.585 2244.530 69.415 ;
        RECT 5.330 61.145 2244.530 63.975 ;
        RECT 5.330 55.705 2244.530 58.535 ;
        RECT 5.330 50.265 2244.530 53.095 ;
        RECT 5.330 44.825 2244.530 47.655 ;
        RECT 5.330 39.385 2244.530 42.215 ;
        RECT 5.330 33.945 2244.530 36.775 ;
        RECT 5.330 28.505 2244.530 31.335 ;
        RECT 5.330 23.065 2244.530 25.895 ;
        RECT 5.330 17.625 2244.530 20.455 ;
        RECT 5.330 12.185 2244.530 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 2244.340 2238.645 ;
      LAYER met1 ;
        RECT 5.520 9.900 2244.340 2238.800 ;
      LAYER met2 ;
        RECT 7.920 4.280 2173.010 2238.745 ;
        RECT 7.920 4.000 106.070 4.280 ;
        RECT 106.910 4.000 110.210 4.280 ;
        RECT 111.050 4.000 114.350 4.280 ;
        RECT 115.190 4.000 118.490 4.280 ;
        RECT 119.330 4.000 122.630 4.280 ;
        RECT 123.470 4.000 126.770 4.280 ;
        RECT 127.610 4.000 130.910 4.280 ;
        RECT 131.750 4.000 135.050 4.280 ;
        RECT 135.890 4.000 139.190 4.280 ;
        RECT 140.030 4.000 143.330 4.280 ;
        RECT 144.170 4.000 147.470 4.280 ;
        RECT 148.310 4.000 151.610 4.280 ;
        RECT 152.450 4.000 155.750 4.280 ;
        RECT 156.590 4.000 159.890 4.280 ;
        RECT 160.730 4.000 164.030 4.280 ;
        RECT 164.870 4.000 168.170 4.280 ;
        RECT 169.010 4.000 172.310 4.280 ;
        RECT 173.150 4.000 176.450 4.280 ;
        RECT 177.290 4.000 180.590 4.280 ;
        RECT 181.430 4.000 184.730 4.280 ;
        RECT 185.570 4.000 188.870 4.280 ;
        RECT 189.710 4.000 193.010 4.280 ;
        RECT 193.850 4.000 197.150 4.280 ;
        RECT 197.990 4.000 201.290 4.280 ;
        RECT 202.130 4.000 205.430 4.280 ;
        RECT 206.270 4.000 209.570 4.280 ;
        RECT 210.410 4.000 213.710 4.280 ;
        RECT 214.550 4.000 217.850 4.280 ;
        RECT 218.690 4.000 221.990 4.280 ;
        RECT 222.830 4.000 226.130 4.280 ;
        RECT 226.970 4.000 230.270 4.280 ;
        RECT 231.110 4.000 234.410 4.280 ;
        RECT 235.250 4.000 238.550 4.280 ;
        RECT 239.390 4.000 242.690 4.280 ;
        RECT 243.530 4.000 246.830 4.280 ;
        RECT 247.670 4.000 250.970 4.280 ;
        RECT 251.810 4.000 255.110 4.280 ;
        RECT 255.950 4.000 259.250 4.280 ;
        RECT 260.090 4.000 263.390 4.280 ;
        RECT 264.230 4.000 267.530 4.280 ;
        RECT 268.370 4.000 271.670 4.280 ;
        RECT 272.510 4.000 275.810 4.280 ;
        RECT 276.650 4.000 279.950 4.280 ;
        RECT 280.790 4.000 284.090 4.280 ;
        RECT 284.930 4.000 288.230 4.280 ;
        RECT 289.070 4.000 292.370 4.280 ;
        RECT 293.210 4.000 296.510 4.280 ;
        RECT 297.350 4.000 300.650 4.280 ;
        RECT 301.490 4.000 304.790 4.280 ;
        RECT 305.630 4.000 308.930 4.280 ;
        RECT 309.770 4.000 313.070 4.280 ;
        RECT 313.910 4.000 317.210 4.280 ;
        RECT 318.050 4.000 321.350 4.280 ;
        RECT 322.190 4.000 325.490 4.280 ;
        RECT 326.330 4.000 329.630 4.280 ;
        RECT 330.470 4.000 333.770 4.280 ;
        RECT 334.610 4.000 337.910 4.280 ;
        RECT 338.750 4.000 342.050 4.280 ;
        RECT 342.890 4.000 346.190 4.280 ;
        RECT 347.030 4.000 350.330 4.280 ;
        RECT 351.170 4.000 354.470 4.280 ;
        RECT 355.310 4.000 358.610 4.280 ;
        RECT 359.450 4.000 362.750 4.280 ;
        RECT 363.590 4.000 366.890 4.280 ;
        RECT 367.730 4.000 371.030 4.280 ;
        RECT 371.870 4.000 375.170 4.280 ;
        RECT 376.010 4.000 379.310 4.280 ;
        RECT 380.150 4.000 383.450 4.280 ;
        RECT 384.290 4.000 387.590 4.280 ;
        RECT 388.430 4.000 391.730 4.280 ;
        RECT 392.570 4.000 395.870 4.280 ;
        RECT 396.710 4.000 400.010 4.280 ;
        RECT 400.850 4.000 404.150 4.280 ;
        RECT 404.990 4.000 408.290 4.280 ;
        RECT 409.130 4.000 412.430 4.280 ;
        RECT 413.270 4.000 416.570 4.280 ;
        RECT 417.410 4.000 420.710 4.280 ;
        RECT 421.550 4.000 424.850 4.280 ;
        RECT 425.690 4.000 428.990 4.280 ;
        RECT 429.830 4.000 433.130 4.280 ;
        RECT 433.970 4.000 437.270 4.280 ;
        RECT 438.110 4.000 441.410 4.280 ;
        RECT 442.250 4.000 445.550 4.280 ;
        RECT 446.390 4.000 449.690 4.280 ;
        RECT 450.530 4.000 453.830 4.280 ;
        RECT 454.670 4.000 457.970 4.280 ;
        RECT 458.810 4.000 462.110 4.280 ;
        RECT 462.950 4.000 466.250 4.280 ;
        RECT 467.090 4.000 470.390 4.280 ;
        RECT 471.230 4.000 474.530 4.280 ;
        RECT 475.370 4.000 478.670 4.280 ;
        RECT 479.510 4.000 482.810 4.280 ;
        RECT 483.650 4.000 486.950 4.280 ;
        RECT 487.790 4.000 491.090 4.280 ;
        RECT 491.930 4.000 495.230 4.280 ;
        RECT 496.070 4.000 499.370 4.280 ;
        RECT 500.210 4.000 503.510 4.280 ;
        RECT 504.350 4.000 507.650 4.280 ;
        RECT 508.490 4.000 511.790 4.280 ;
        RECT 512.630 4.000 515.930 4.280 ;
        RECT 516.770 4.000 520.070 4.280 ;
        RECT 520.910 4.000 524.210 4.280 ;
        RECT 525.050 4.000 528.350 4.280 ;
        RECT 529.190 4.000 532.490 4.280 ;
        RECT 533.330 4.000 536.630 4.280 ;
        RECT 537.470 4.000 540.770 4.280 ;
        RECT 541.610 4.000 544.910 4.280 ;
        RECT 545.750 4.000 549.050 4.280 ;
        RECT 549.890 4.000 553.190 4.280 ;
        RECT 554.030 4.000 557.330 4.280 ;
        RECT 558.170 4.000 561.470 4.280 ;
        RECT 562.310 4.000 565.610 4.280 ;
        RECT 566.450 4.000 569.750 4.280 ;
        RECT 570.590 4.000 573.890 4.280 ;
        RECT 574.730 4.000 578.030 4.280 ;
        RECT 578.870 4.000 582.170 4.280 ;
        RECT 583.010 4.000 586.310 4.280 ;
        RECT 587.150 4.000 590.450 4.280 ;
        RECT 591.290 4.000 594.590 4.280 ;
        RECT 595.430 4.000 598.730 4.280 ;
        RECT 599.570 4.000 602.870 4.280 ;
        RECT 603.710 4.000 607.010 4.280 ;
        RECT 607.850 4.000 611.150 4.280 ;
        RECT 611.990 4.000 615.290 4.280 ;
        RECT 616.130 4.000 619.430 4.280 ;
        RECT 620.270 4.000 623.570 4.280 ;
        RECT 624.410 4.000 627.710 4.280 ;
        RECT 628.550 4.000 631.850 4.280 ;
        RECT 632.690 4.000 635.990 4.280 ;
        RECT 636.830 4.000 640.130 4.280 ;
        RECT 640.970 4.000 644.270 4.280 ;
        RECT 645.110 4.000 648.410 4.280 ;
        RECT 649.250 4.000 652.550 4.280 ;
        RECT 653.390 4.000 656.690 4.280 ;
        RECT 657.530 4.000 660.830 4.280 ;
        RECT 661.670 4.000 664.970 4.280 ;
        RECT 665.810 4.000 669.110 4.280 ;
        RECT 669.950 4.000 673.250 4.280 ;
        RECT 674.090 4.000 677.390 4.280 ;
        RECT 678.230 4.000 681.530 4.280 ;
        RECT 682.370 4.000 685.670 4.280 ;
        RECT 686.510 4.000 689.810 4.280 ;
        RECT 690.650 4.000 693.950 4.280 ;
        RECT 694.790 4.000 698.090 4.280 ;
        RECT 698.930 4.000 702.230 4.280 ;
        RECT 703.070 4.000 706.370 4.280 ;
        RECT 707.210 4.000 710.510 4.280 ;
        RECT 711.350 4.000 714.650 4.280 ;
        RECT 715.490 4.000 718.790 4.280 ;
        RECT 719.630 4.000 722.930 4.280 ;
        RECT 723.770 4.000 727.070 4.280 ;
        RECT 727.910 4.000 731.210 4.280 ;
        RECT 732.050 4.000 735.350 4.280 ;
        RECT 736.190 4.000 739.490 4.280 ;
        RECT 740.330 4.000 743.630 4.280 ;
        RECT 744.470 4.000 747.770 4.280 ;
        RECT 748.610 4.000 751.910 4.280 ;
        RECT 752.750 4.000 756.050 4.280 ;
        RECT 756.890 4.000 760.190 4.280 ;
        RECT 761.030 4.000 764.330 4.280 ;
        RECT 765.170 4.000 768.470 4.280 ;
        RECT 769.310 4.000 772.610 4.280 ;
        RECT 773.450 4.000 776.750 4.280 ;
        RECT 777.590 4.000 780.890 4.280 ;
        RECT 781.730 4.000 785.030 4.280 ;
        RECT 785.870 4.000 789.170 4.280 ;
        RECT 790.010 4.000 793.310 4.280 ;
        RECT 794.150 4.000 797.450 4.280 ;
        RECT 798.290 4.000 801.590 4.280 ;
        RECT 802.430 4.000 805.730 4.280 ;
        RECT 806.570 4.000 809.870 4.280 ;
        RECT 810.710 4.000 814.010 4.280 ;
        RECT 814.850 4.000 818.150 4.280 ;
        RECT 818.990 4.000 822.290 4.280 ;
        RECT 823.130 4.000 826.430 4.280 ;
        RECT 827.270 4.000 830.570 4.280 ;
        RECT 831.410 4.000 834.710 4.280 ;
        RECT 835.550 4.000 838.850 4.280 ;
        RECT 839.690 4.000 842.990 4.280 ;
        RECT 843.830 4.000 847.130 4.280 ;
        RECT 847.970 4.000 851.270 4.280 ;
        RECT 852.110 4.000 855.410 4.280 ;
        RECT 856.250 4.000 859.550 4.280 ;
        RECT 860.390 4.000 863.690 4.280 ;
        RECT 864.530 4.000 867.830 4.280 ;
        RECT 868.670 4.000 871.970 4.280 ;
        RECT 872.810 4.000 876.110 4.280 ;
        RECT 876.950 4.000 880.250 4.280 ;
        RECT 881.090 4.000 884.390 4.280 ;
        RECT 885.230 4.000 888.530 4.280 ;
        RECT 889.370 4.000 892.670 4.280 ;
        RECT 893.510 4.000 896.810 4.280 ;
        RECT 897.650 4.000 900.950 4.280 ;
        RECT 901.790 4.000 905.090 4.280 ;
        RECT 905.930 4.000 909.230 4.280 ;
        RECT 910.070 4.000 913.370 4.280 ;
        RECT 914.210 4.000 917.510 4.280 ;
        RECT 918.350 4.000 921.650 4.280 ;
        RECT 922.490 4.000 925.790 4.280 ;
        RECT 926.630 4.000 929.930 4.280 ;
        RECT 930.770 4.000 934.070 4.280 ;
        RECT 934.910 4.000 938.210 4.280 ;
        RECT 939.050 4.000 942.350 4.280 ;
        RECT 943.190 4.000 946.490 4.280 ;
        RECT 947.330 4.000 950.630 4.280 ;
        RECT 951.470 4.000 954.770 4.280 ;
        RECT 955.610 4.000 958.910 4.280 ;
        RECT 959.750 4.000 963.050 4.280 ;
        RECT 963.890 4.000 967.190 4.280 ;
        RECT 968.030 4.000 971.330 4.280 ;
        RECT 972.170 4.000 975.470 4.280 ;
        RECT 976.310 4.000 979.610 4.280 ;
        RECT 980.450 4.000 983.750 4.280 ;
        RECT 984.590 4.000 987.890 4.280 ;
        RECT 988.730 4.000 992.030 4.280 ;
        RECT 992.870 4.000 996.170 4.280 ;
        RECT 997.010 4.000 1000.310 4.280 ;
        RECT 1001.150 4.000 1004.450 4.280 ;
        RECT 1005.290 4.000 1008.590 4.280 ;
        RECT 1009.430 4.000 1012.730 4.280 ;
        RECT 1013.570 4.000 1016.870 4.280 ;
        RECT 1017.710 4.000 1021.010 4.280 ;
        RECT 1021.850 4.000 1025.150 4.280 ;
        RECT 1025.990 4.000 1029.290 4.280 ;
        RECT 1030.130 4.000 1033.430 4.280 ;
        RECT 1034.270 4.000 1037.570 4.280 ;
        RECT 1038.410 4.000 1041.710 4.280 ;
        RECT 1042.550 4.000 1045.850 4.280 ;
        RECT 1046.690 4.000 1049.990 4.280 ;
        RECT 1050.830 4.000 1054.130 4.280 ;
        RECT 1054.970 4.000 1058.270 4.280 ;
        RECT 1059.110 4.000 1062.410 4.280 ;
        RECT 1063.250 4.000 1066.550 4.280 ;
        RECT 1067.390 4.000 1070.690 4.280 ;
        RECT 1071.530 4.000 1074.830 4.280 ;
        RECT 1075.670 4.000 1078.970 4.280 ;
        RECT 1079.810 4.000 1083.110 4.280 ;
        RECT 1083.950 4.000 1087.250 4.280 ;
        RECT 1088.090 4.000 1091.390 4.280 ;
        RECT 1092.230 4.000 1095.530 4.280 ;
        RECT 1096.370 4.000 1099.670 4.280 ;
        RECT 1100.510 4.000 1103.810 4.280 ;
        RECT 1104.650 4.000 1107.950 4.280 ;
        RECT 1108.790 4.000 1112.090 4.280 ;
        RECT 1112.930 4.000 1116.230 4.280 ;
        RECT 1117.070 4.000 1120.370 4.280 ;
        RECT 1121.210 4.000 1124.510 4.280 ;
        RECT 1125.350 4.000 1128.650 4.280 ;
        RECT 1129.490 4.000 1132.790 4.280 ;
        RECT 1133.630 4.000 1136.930 4.280 ;
        RECT 1137.770 4.000 1141.070 4.280 ;
        RECT 1141.910 4.000 1145.210 4.280 ;
        RECT 1146.050 4.000 1149.350 4.280 ;
        RECT 1150.190 4.000 1153.490 4.280 ;
        RECT 1154.330 4.000 1157.630 4.280 ;
        RECT 1158.470 4.000 1161.770 4.280 ;
        RECT 1162.610 4.000 1165.910 4.280 ;
        RECT 1166.750 4.000 1170.050 4.280 ;
        RECT 1170.890 4.000 1174.190 4.280 ;
        RECT 1175.030 4.000 1178.330 4.280 ;
        RECT 1179.170 4.000 1182.470 4.280 ;
        RECT 1183.310 4.000 1186.610 4.280 ;
        RECT 1187.450 4.000 1190.750 4.280 ;
        RECT 1191.590 4.000 1194.890 4.280 ;
        RECT 1195.730 4.000 1199.030 4.280 ;
        RECT 1199.870 4.000 1203.170 4.280 ;
        RECT 1204.010 4.000 1207.310 4.280 ;
        RECT 1208.150 4.000 1211.450 4.280 ;
        RECT 1212.290 4.000 1215.590 4.280 ;
        RECT 1216.430 4.000 1219.730 4.280 ;
        RECT 1220.570 4.000 1223.870 4.280 ;
        RECT 1224.710 4.000 1228.010 4.280 ;
        RECT 1228.850 4.000 1232.150 4.280 ;
        RECT 1232.990 4.000 1236.290 4.280 ;
        RECT 1237.130 4.000 1240.430 4.280 ;
        RECT 1241.270 4.000 1244.570 4.280 ;
        RECT 1245.410 4.000 1248.710 4.280 ;
        RECT 1249.550 4.000 1252.850 4.280 ;
        RECT 1253.690 4.000 1256.990 4.280 ;
        RECT 1257.830 4.000 1261.130 4.280 ;
        RECT 1261.970 4.000 1265.270 4.280 ;
        RECT 1266.110 4.000 1269.410 4.280 ;
        RECT 1270.250 4.000 1273.550 4.280 ;
        RECT 1274.390 4.000 1277.690 4.280 ;
        RECT 1278.530 4.000 1281.830 4.280 ;
        RECT 1282.670 4.000 1285.970 4.280 ;
        RECT 1286.810 4.000 1290.110 4.280 ;
        RECT 1290.950 4.000 1294.250 4.280 ;
        RECT 1295.090 4.000 1298.390 4.280 ;
        RECT 1299.230 4.000 1302.530 4.280 ;
        RECT 1303.370 4.000 1306.670 4.280 ;
        RECT 1307.510 4.000 1310.810 4.280 ;
        RECT 1311.650 4.000 1314.950 4.280 ;
        RECT 1315.790 4.000 1319.090 4.280 ;
        RECT 1319.930 4.000 1323.230 4.280 ;
        RECT 1324.070 4.000 1327.370 4.280 ;
        RECT 1328.210 4.000 1331.510 4.280 ;
        RECT 1332.350 4.000 1335.650 4.280 ;
        RECT 1336.490 4.000 1339.790 4.280 ;
        RECT 1340.630 4.000 1343.930 4.280 ;
        RECT 1344.770 4.000 1348.070 4.280 ;
        RECT 1348.910 4.000 1352.210 4.280 ;
        RECT 1353.050 4.000 1356.350 4.280 ;
        RECT 1357.190 4.000 1360.490 4.280 ;
        RECT 1361.330 4.000 1364.630 4.280 ;
        RECT 1365.470 4.000 1368.770 4.280 ;
        RECT 1369.610 4.000 1372.910 4.280 ;
        RECT 1373.750 4.000 1377.050 4.280 ;
        RECT 1377.890 4.000 1381.190 4.280 ;
        RECT 1382.030 4.000 1385.330 4.280 ;
        RECT 1386.170 4.000 1389.470 4.280 ;
        RECT 1390.310 4.000 1393.610 4.280 ;
        RECT 1394.450 4.000 1397.750 4.280 ;
        RECT 1398.590 4.000 1401.890 4.280 ;
        RECT 1402.730 4.000 1406.030 4.280 ;
        RECT 1406.870 4.000 1410.170 4.280 ;
        RECT 1411.010 4.000 1414.310 4.280 ;
        RECT 1415.150 4.000 1418.450 4.280 ;
        RECT 1419.290 4.000 1422.590 4.280 ;
        RECT 1423.430 4.000 1426.730 4.280 ;
        RECT 1427.570 4.000 1430.870 4.280 ;
        RECT 1431.710 4.000 1435.010 4.280 ;
        RECT 1435.850 4.000 1439.150 4.280 ;
        RECT 1439.990 4.000 1443.290 4.280 ;
        RECT 1444.130 4.000 1447.430 4.280 ;
        RECT 1448.270 4.000 1451.570 4.280 ;
        RECT 1452.410 4.000 1455.710 4.280 ;
        RECT 1456.550 4.000 1459.850 4.280 ;
        RECT 1460.690 4.000 1463.990 4.280 ;
        RECT 1464.830 4.000 1468.130 4.280 ;
        RECT 1468.970 4.000 1472.270 4.280 ;
        RECT 1473.110 4.000 1476.410 4.280 ;
        RECT 1477.250 4.000 1480.550 4.280 ;
        RECT 1481.390 4.000 1484.690 4.280 ;
        RECT 1485.530 4.000 1488.830 4.280 ;
        RECT 1489.670 4.000 1492.970 4.280 ;
        RECT 1493.810 4.000 1497.110 4.280 ;
        RECT 1497.950 4.000 1501.250 4.280 ;
        RECT 1502.090 4.000 1505.390 4.280 ;
        RECT 1506.230 4.000 1509.530 4.280 ;
        RECT 1510.370 4.000 1513.670 4.280 ;
        RECT 1514.510 4.000 1517.810 4.280 ;
        RECT 1518.650 4.000 1521.950 4.280 ;
        RECT 1522.790 4.000 1526.090 4.280 ;
        RECT 1526.930 4.000 1530.230 4.280 ;
        RECT 1531.070 4.000 1534.370 4.280 ;
        RECT 1535.210 4.000 1538.510 4.280 ;
        RECT 1539.350 4.000 1542.650 4.280 ;
        RECT 1543.490 4.000 1546.790 4.280 ;
        RECT 1547.630 4.000 1550.930 4.280 ;
        RECT 1551.770 4.000 1555.070 4.280 ;
        RECT 1555.910 4.000 1559.210 4.280 ;
        RECT 1560.050 4.000 1563.350 4.280 ;
        RECT 1564.190 4.000 1567.490 4.280 ;
        RECT 1568.330 4.000 1571.630 4.280 ;
        RECT 1572.470 4.000 1575.770 4.280 ;
        RECT 1576.610 4.000 1579.910 4.280 ;
        RECT 1580.750 4.000 1584.050 4.280 ;
        RECT 1584.890 4.000 1588.190 4.280 ;
        RECT 1589.030 4.000 1592.330 4.280 ;
        RECT 1593.170 4.000 1596.470 4.280 ;
        RECT 1597.310 4.000 1600.610 4.280 ;
        RECT 1601.450 4.000 1604.750 4.280 ;
        RECT 1605.590 4.000 1608.890 4.280 ;
        RECT 1609.730 4.000 1613.030 4.280 ;
        RECT 1613.870 4.000 1617.170 4.280 ;
        RECT 1618.010 4.000 1621.310 4.280 ;
        RECT 1622.150 4.000 1625.450 4.280 ;
        RECT 1626.290 4.000 1629.590 4.280 ;
        RECT 1630.430 4.000 1633.730 4.280 ;
        RECT 1634.570 4.000 1637.870 4.280 ;
        RECT 1638.710 4.000 1642.010 4.280 ;
        RECT 1642.850 4.000 1646.150 4.280 ;
        RECT 1646.990 4.000 1650.290 4.280 ;
        RECT 1651.130 4.000 1654.430 4.280 ;
        RECT 1655.270 4.000 1658.570 4.280 ;
        RECT 1659.410 4.000 1662.710 4.280 ;
        RECT 1663.550 4.000 1666.850 4.280 ;
        RECT 1667.690 4.000 1670.990 4.280 ;
        RECT 1671.830 4.000 1675.130 4.280 ;
        RECT 1675.970 4.000 1679.270 4.280 ;
        RECT 1680.110 4.000 1683.410 4.280 ;
        RECT 1684.250 4.000 1687.550 4.280 ;
        RECT 1688.390 4.000 1691.690 4.280 ;
        RECT 1692.530 4.000 1695.830 4.280 ;
        RECT 1696.670 4.000 1699.970 4.280 ;
        RECT 1700.810 4.000 1704.110 4.280 ;
        RECT 1704.950 4.000 1708.250 4.280 ;
        RECT 1709.090 4.000 1712.390 4.280 ;
        RECT 1713.230 4.000 1716.530 4.280 ;
        RECT 1717.370 4.000 1720.670 4.280 ;
        RECT 1721.510 4.000 1724.810 4.280 ;
        RECT 1725.650 4.000 1728.950 4.280 ;
        RECT 1729.790 4.000 1733.090 4.280 ;
        RECT 1733.930 4.000 1737.230 4.280 ;
        RECT 1738.070 4.000 1741.370 4.280 ;
        RECT 1742.210 4.000 1745.510 4.280 ;
        RECT 1746.350 4.000 1749.650 4.280 ;
        RECT 1750.490 4.000 1753.790 4.280 ;
        RECT 1754.630 4.000 1757.930 4.280 ;
        RECT 1758.770 4.000 1762.070 4.280 ;
        RECT 1762.910 4.000 1766.210 4.280 ;
        RECT 1767.050 4.000 1770.350 4.280 ;
        RECT 1771.190 4.000 1774.490 4.280 ;
        RECT 1775.330 4.000 1778.630 4.280 ;
        RECT 1779.470 4.000 1782.770 4.280 ;
        RECT 1783.610 4.000 1786.910 4.280 ;
        RECT 1787.750 4.000 1791.050 4.280 ;
        RECT 1791.890 4.000 1795.190 4.280 ;
        RECT 1796.030 4.000 1799.330 4.280 ;
        RECT 1800.170 4.000 1803.470 4.280 ;
        RECT 1804.310 4.000 1807.610 4.280 ;
        RECT 1808.450 4.000 1811.750 4.280 ;
        RECT 1812.590 4.000 1815.890 4.280 ;
        RECT 1816.730 4.000 1820.030 4.280 ;
        RECT 1820.870 4.000 1824.170 4.280 ;
        RECT 1825.010 4.000 1828.310 4.280 ;
        RECT 1829.150 4.000 1832.450 4.280 ;
        RECT 1833.290 4.000 1836.590 4.280 ;
        RECT 1837.430 4.000 1840.730 4.280 ;
        RECT 1841.570 4.000 1844.870 4.280 ;
        RECT 1845.710 4.000 1849.010 4.280 ;
        RECT 1849.850 4.000 1853.150 4.280 ;
        RECT 1853.990 4.000 1857.290 4.280 ;
        RECT 1858.130 4.000 1861.430 4.280 ;
        RECT 1862.270 4.000 1865.570 4.280 ;
        RECT 1866.410 4.000 1869.710 4.280 ;
        RECT 1870.550 4.000 1873.850 4.280 ;
        RECT 1874.690 4.000 1877.990 4.280 ;
        RECT 1878.830 4.000 1882.130 4.280 ;
        RECT 1882.970 4.000 1886.270 4.280 ;
        RECT 1887.110 4.000 1890.410 4.280 ;
        RECT 1891.250 4.000 1894.550 4.280 ;
        RECT 1895.390 4.000 1898.690 4.280 ;
        RECT 1899.530 4.000 1902.830 4.280 ;
        RECT 1903.670 4.000 1906.970 4.280 ;
        RECT 1907.810 4.000 1911.110 4.280 ;
        RECT 1911.950 4.000 1915.250 4.280 ;
        RECT 1916.090 4.000 1919.390 4.280 ;
        RECT 1920.230 4.000 1923.530 4.280 ;
        RECT 1924.370 4.000 1927.670 4.280 ;
        RECT 1928.510 4.000 1931.810 4.280 ;
        RECT 1932.650 4.000 1935.950 4.280 ;
        RECT 1936.790 4.000 1940.090 4.280 ;
        RECT 1940.930 4.000 1944.230 4.280 ;
        RECT 1945.070 4.000 1948.370 4.280 ;
        RECT 1949.210 4.000 1952.510 4.280 ;
        RECT 1953.350 4.000 1956.650 4.280 ;
        RECT 1957.490 4.000 1960.790 4.280 ;
        RECT 1961.630 4.000 1964.930 4.280 ;
        RECT 1965.770 4.000 1969.070 4.280 ;
        RECT 1969.910 4.000 1973.210 4.280 ;
        RECT 1974.050 4.000 1977.350 4.280 ;
        RECT 1978.190 4.000 1981.490 4.280 ;
        RECT 1982.330 4.000 1985.630 4.280 ;
        RECT 1986.470 4.000 1989.770 4.280 ;
        RECT 1990.610 4.000 1993.910 4.280 ;
        RECT 1994.750 4.000 1998.050 4.280 ;
        RECT 1998.890 4.000 2002.190 4.280 ;
        RECT 2003.030 4.000 2006.330 4.280 ;
        RECT 2007.170 4.000 2010.470 4.280 ;
        RECT 2011.310 4.000 2014.610 4.280 ;
        RECT 2015.450 4.000 2018.750 4.280 ;
        RECT 2019.590 4.000 2022.890 4.280 ;
        RECT 2023.730 4.000 2027.030 4.280 ;
        RECT 2027.870 4.000 2031.170 4.280 ;
        RECT 2032.010 4.000 2035.310 4.280 ;
        RECT 2036.150 4.000 2039.450 4.280 ;
        RECT 2040.290 4.000 2043.590 4.280 ;
        RECT 2044.430 4.000 2047.730 4.280 ;
        RECT 2048.570 4.000 2051.870 4.280 ;
        RECT 2052.710 4.000 2056.010 4.280 ;
        RECT 2056.850 4.000 2060.150 4.280 ;
        RECT 2060.990 4.000 2064.290 4.280 ;
        RECT 2065.130 4.000 2068.430 4.280 ;
        RECT 2069.270 4.000 2072.570 4.280 ;
        RECT 2073.410 4.000 2076.710 4.280 ;
        RECT 2077.550 4.000 2080.850 4.280 ;
        RECT 2081.690 4.000 2084.990 4.280 ;
        RECT 2085.830 4.000 2089.130 4.280 ;
        RECT 2089.970 4.000 2093.270 4.280 ;
        RECT 2094.110 4.000 2097.410 4.280 ;
        RECT 2098.250 4.000 2101.550 4.280 ;
        RECT 2102.390 4.000 2105.690 4.280 ;
        RECT 2106.530 4.000 2109.830 4.280 ;
        RECT 2110.670 4.000 2113.970 4.280 ;
        RECT 2114.810 4.000 2118.110 4.280 ;
        RECT 2118.950 4.000 2122.250 4.280 ;
        RECT 2123.090 4.000 2126.390 4.280 ;
        RECT 2127.230 4.000 2130.530 4.280 ;
        RECT 2131.370 4.000 2134.670 4.280 ;
        RECT 2135.510 4.000 2138.810 4.280 ;
        RECT 2139.650 4.000 2142.950 4.280 ;
        RECT 2143.790 4.000 2173.010 4.280 ;
      LAYER met3 ;
        RECT 21.050 10.715 2173.030 2238.725 ;
      LAYER met4 ;
        RECT 278.135 44.375 327.840 721.305 ;
        RECT 330.240 44.375 404.640 721.305 ;
        RECT 407.040 44.375 481.440 721.305 ;
        RECT 483.840 44.375 558.240 721.305 ;
        RECT 560.640 44.375 635.040 721.305 ;
        RECT 637.440 44.375 640.025 721.305 ;
  END
END user_proj_example
END LIBRARY

