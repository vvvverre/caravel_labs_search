// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module user_proj_example #(
    parameter SEQ_WIDTH = 72,
    parameter E_WIDTH = 20,

    parameter STAGE_WIDTH = 8,
    parameter PARALLEL_UNITS = 1
)(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IRQ
    output [2:0] irq
);
    wire clk;
    wire rst;

    // IRQ
    assign irq = 3'b000;	// Unused

    // LA
    // assign la_data_out = {{(127-BITS){1'b0}}, count};
    // Assuming LA probes [63:32] are for controlling the count register  
    // assign la_write = ~la_oenb[63:32] & ~{BITS{valid}};
    // Assuming LA probes [65:64] are for controlling the count clk & reset  
    assign clk = wb_clk_i;
    assign rst = wb_rst_i;


    wb_find #
    (
        .SEQ_WIDTH(SEQ_WIDTH),
        .E_WIDTH(E_WIDTH),

        .STAGE_WIDTH(STAGE_WIDTH),
        .PARALLEL_UNITS(PARALLEL_UNITS)
    ) inst_wb_find (
        .wb_clk_i(clk),
        .wb_rst_i(rst),

        .wbs_stb_i(wbs_stb_i),
        .wbs_cyc_i(wbs_cyc_i),

        .wbs_we_i(wbs_we_i),
        .wbs_sel_i(wbs_sel_i),

        .wbs_dat_i(wbs_dat_i),
        .wbs_adr_i(wbs_adr_i),

        .wbs_ack_o(wbs_ack_o),
        .wbs_dat_o(wbs_dat_o),

        .la_data_in(la_data_in),
        .la_data_out(la_data_out),
        .la_oenb(la_oenb)
    );
    

endmodule
`default_nettype wire
